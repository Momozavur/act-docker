magic
tech scmos
timestamp 1761015633
<< nwell >>
rect -11 -1 74 51
<< pwell >>
rect -11 52 74 81
rect -11 -25 74 -2
<< ntransistor >>
rect 10 58 12 63
rect 16 58 18 63
rect 26 58 28 63
rect 33 58 35 63
rect 51 58 53 63
rect 60 58 62 63
rect 10 -13 12 -8
rect 19 -13 21 -8
rect 37 -13 39 -8
rect 43 -13 45 -8
rect 52 -13 54 -8
rect 58 -13 60 -8
<< ptransistor >>
rect 10 35 12 45
rect 16 35 18 45
rect 26 35 28 45
rect 33 35 35 45
rect 51 35 53 45
rect 60 35 62 45
rect 10 5 12 15
rect 19 5 21 15
rect 37 5 39 15
rect 43 5 45 15
rect 52 5 54 15
rect 58 5 60 15
<< ndiffusion >>
rect 9 58 10 63
rect 12 58 16 63
rect 18 58 19 63
rect 25 58 26 63
rect 28 58 33 63
rect 35 58 36 63
rect 50 58 51 63
rect 53 58 54 63
rect 59 58 60 63
rect 62 58 63 63
rect 9 -13 10 -8
rect 12 -13 13 -8
rect 18 -13 19 -8
rect 21 -13 22 -8
rect 36 -13 37 -8
rect 39 -13 43 -8
rect 45 -13 46 -8
rect 51 -13 52 -8
rect 54 -13 58 -8
rect 60 -13 61 -8
<< pdiffusion >>
rect 9 35 10 45
rect 12 35 16 45
rect 18 35 19 45
rect 25 35 26 45
rect 28 35 33 45
rect 35 35 36 45
rect 50 35 51 45
rect 53 35 54 45
rect 59 35 60 45
rect 62 35 63 45
rect 9 5 10 15
rect 12 5 13 15
rect 18 5 19 15
rect 21 5 22 15
rect 36 5 37 15
rect 39 5 43 15
rect 45 5 46 15
rect 51 5 52 15
rect 54 5 58 15
rect 60 5 61 15
<< ndcontact >>
rect 19 58 25 63
rect 45 58 50 63
rect 63 58 68 63
rect 4 -13 9 -8
rect 22 -13 27 -8
rect 31 -13 36 -8
rect 61 -13 66 -8
<< pdcontact >>
rect 19 35 25 45
rect 45 35 50 45
rect 63 35 68 45
rect 4 5 9 15
rect 22 5 27 15
rect 31 5 36 15
rect 61 5 66 15
<< psubstratepcontact >>
rect 1 67 13 72
rect 1 -22 9 -17
<< nsubstratencontact >>
rect 1 26 13 31
rect 42 19 51 24
<< polysilicon >>
rect 51 75 68 77
rect 16 69 42 71
rect 10 63 12 66
rect 16 63 18 69
rect 40 67 42 69
rect 51 67 53 75
rect 26 63 28 66
rect 33 63 35 66
rect 40 65 53 67
rect 66 66 68 75
rect 51 63 53 65
rect 60 63 62 66
rect 10 45 12 58
rect 16 55 18 58
rect 26 57 28 58
rect 21 55 28 57
rect 21 48 23 55
rect 33 54 35 58
rect 16 46 23 48
rect 16 45 18 46
rect 26 45 28 48
rect 33 45 35 49
rect 51 45 53 58
rect 60 45 62 58
rect 10 32 12 35
rect 16 32 18 35
rect 26 29 28 35
rect 33 32 35 35
rect 51 34 53 35
rect 47 32 53 34
rect 47 29 49 32
rect 60 29 62 35
rect 26 27 49 29
rect 52 27 62 29
rect 1 21 21 23
rect 10 15 12 18
rect 19 15 21 21
rect 37 15 39 18
rect 43 15 45 18
rect 52 15 54 27
rect 58 15 60 18
rect 10 -8 12 5
rect 19 -8 21 5
rect 37 2 39 5
rect 43 4 45 5
rect 52 4 54 5
rect 43 2 54 4
rect 58 2 60 5
rect 37 -8 39 -5
rect 43 -8 45 2
rect 52 -8 54 2
rect 58 -8 60 -5
rect 10 -14 12 -13
rect -6 -16 12 -14
rect 19 -14 21 -13
rect 37 -14 39 -13
rect 19 -16 39 -14
rect 43 -16 45 -13
rect 52 -16 54 -13
rect 10 -19 12 -16
rect 58 -19 60 -13
rect 10 -21 60 -19
<< polycontact >>
rect 57 66 62 71
rect 68 66 73 71
rect 5 49 10 54
rect 16 27 21 32
rect -4 18 1 23
rect 34 18 39 23
rect -11 -19 -6 -14
<< metal1 >>
rect 4 63 9 67
rect 19 66 57 71
rect 19 63 25 66
rect -11 49 5 54
rect 19 45 25 58
rect 45 45 50 58
rect 63 54 68 58
rect 59 49 68 54
rect 63 45 68 49
rect 4 31 9 35
rect 45 32 50 35
rect 21 27 50 32
rect 4 23 9 26
rect 9 18 18 23
rect 0 13 1 18
rect 13 15 18 18
rect 22 18 34 23
rect 22 15 27 18
rect 46 15 51 19
rect 4 1 9 5
rect 4 -8 9 -4
rect 22 -8 27 5
rect 31 -8 36 5
rect 61 -3 66 5
rect 61 -8 74 -3
rect 69 -13 74 -8
rect 13 -17 18 -13
rect 31 -17 36 -13
rect 9 -22 22 -17
rect 72 -22 74 -17
<< m2contact >>
rect 54 49 59 54
rect 4 -4 9 1
rect -11 -24 -6 -19
rect 31 -22 36 -17
rect 67 -22 72 -17
<< pm12contact >>
rect 33 49 38 54
rect 58 18 63 23
<< pdm12contact >>
rect 4 35 9 45
rect 36 35 41 45
rect 54 35 59 45
rect 13 5 18 15
rect 46 5 51 15
<< ndm12contact >>
rect 4 58 9 63
rect 36 58 41 63
rect 54 58 59 63
rect 13 -13 18 -8
rect 46 -13 51 -8
<< metal2 >>
rect 9 58 36 63
rect 41 58 54 63
rect 59 58 72 63
rect 38 49 54 54
rect 9 35 36 45
rect 41 35 54 45
rect 18 5 46 15
rect 58 1 63 18
rect 9 -4 63 1
rect 67 -8 72 58
rect 18 -13 46 -8
rect 51 -13 72 -8
rect 56 -20 67 -17
rect 36 -22 67 -20
rect 31 -25 61 -22
<< m123contact >>
rect 68 71 73 76
rect 4 18 9 23
rect -5 13 0 18
rect 22 -22 27 -17
<< labels >>
rlabel polysilicon 11 51 11 51 5 in
rlabel polysilicon 11 -2 11 -2 1 r0
rlabel polysilicon 20 -2 20 -2 1 r1
rlabel polysilicon 17 70 17 70 5 w
rlabel psubstratepcontact 7 69 7 69 1 GND!
rlabel nsubstratencontact 6 28 6 28 1 Vdd!
rlabel metal1 63 -6 63 -6 1 port0
rlabel metal1 34 -6 34 -6 1 port1
rlabel metal1 56 68 56 68 1 tmp
<< end >>
