magic
tech scmos
timestamp 1765690562
<< nwell >>
rect 68 53 115 82
<< pwell >>
rect 68 29 115 52
<< ntransistor >>
rect 85 41 87 46
rect 96 41 98 46
<< ptransistor >>
rect 85 60 87 70
rect 96 60 98 70
<< ndiffusion >>
rect 79 41 85 46
rect 87 41 96 46
rect 98 41 104 46
<< pdiffusion >>
rect 79 60 85 70
rect 87 60 89 70
rect 94 60 96 70
rect 98 60 104 70
<< ndcontact >>
rect 74 41 79 46
rect 104 41 109 46
<< pdcontact >>
rect 74 60 79 70
rect 89 60 94 70
rect 104 60 109 70
<< psubstratepcontact >>
rect 89 32 94 37
<< nsubstratencontact >>
rect 89 74 94 79
<< polysilicon >>
rect 85 70 87 73
rect 96 70 98 73
rect 85 46 87 60
rect 96 46 98 60
rect 85 38 87 41
rect 96 38 98 41
<< metal1 >>
rect 74 74 89 79
rect 94 74 115 79
rect 74 70 79 74
rect 104 70 109 74
rect 89 55 94 60
rect 89 50 115 55
rect 104 46 109 50
rect 74 37 79 41
rect 74 32 89 37
rect 94 32 115 37
use inv2  inv2_0
timestamp 1765338958
transform 1 0 118 0 1 42
box -10 -13 20 40
<< labels >>
rlabel metal1 110 74 115 79 7 Vdd!
rlabel polysilicon 85 71 87 73 1 a
<< end >>
