magic
tech scmos
timestamp 1765052771
<< metal1 >>
rect -1 88 141 102
rect 454 94 462 106
rect 804 96 812 108
rect 1154 94 1162 111
rect 1406 97 1414 103
rect 1504 94 1512 103
rect 1756 97 1764 103
rect 1854 96 1862 103
rect 2106 97 2114 103
rect 2204 96 2212 103
rect 2456 97 2464 103
rect 2554 96 2562 103
rect 2806 97 2814 103
rect 2904 96 2912 103
rect 3156 97 3164 103
rect 3254 96 3262 103
rect -1 0 141 48
rect 356 7 361 16
rect 706 7 711 16
rect 1056 7 1061 16
rect 477 0 486 7
rect -207 -142 -195 -134
rect -207 -240 -201 -232
rect 3396 -246 3411 -104
rect 3432 -246 3498 -104
rect 3493 -468 3499 -460
rect -207 -492 -195 -484
rect 3487 -566 3499 -558
rect -207 -590 -201 -582
rect 3493 -818 3499 -810
rect -207 -842 -195 -834
rect 3487 -916 3499 -908
rect -207 -940 -201 -932
rect 3493 -1168 3499 -1160
rect -207 -1192 -195 -1184
rect 3487 -1266 3499 -1258
rect -207 -1290 -201 -1282
rect 3493 -1518 3499 -1510
rect -207 -1542 -195 -1534
rect 3487 -1616 3499 -1608
rect -207 -1640 -201 -1632
rect 3493 -1868 3499 -1860
rect -207 -1892 -195 -1884
rect 3487 -1966 3499 -1958
rect -207 -1990 -201 -1982
rect 3493 -2218 3499 -2210
rect -207 -2242 -196 -2234
rect 3487 -2316 3499 -2308
rect -207 -2340 -201 -2332
rect 3493 -2568 3499 -2560
rect -207 -2592 -195 -2584
rect 3487 -2666 3499 -2658
rect -207 -2690 -201 -2682
rect 3493 -2918 3499 -2910
rect -207 -2942 -195 -2934
rect 3487 -3016 3499 -3008
rect -207 -3040 -201 -3032
rect -206 -3396 -140 -3254
rect -119 -3396 -104 -3254
rect 3493 -3268 3499 -3260
rect 3487 -3366 3499 -3358
rect 3150 -3548 3292 -3500
rect 30 -3603 38 -3591
rect 128 -3603 136 -3597
rect 380 -3603 388 -3591
rect 478 -3603 486 -3597
rect 730 -3603 738 -3591
rect 828 -3603 836 -3597
rect 1080 -3603 1088 -3591
rect 1178 -3603 1186 -3597
rect 1430 -3603 1438 -3591
rect 1528 -3603 1536 -3597
rect 1780 -3603 1788 -3591
rect 1878 -3603 1886 -3597
rect 2130 -3603 2138 -3591
rect 2228 -3603 2236 -3597
rect 2480 -3603 2488 -3591
rect 2578 -3603 2586 -3597
rect 2830 -3603 2838 -3591
rect 2928 -3603 2936 -3597
rect 3150 -3602 3292 -3588
<< m2contact >>
rect -1 48 141 88
rect 3411 -246 3432 -104
rect -140 -3396 -119 -3254
rect 3150 -3588 3292 -3548
<< metal2 >>
rect -192 48 -1 88
rect 141 48 3484 88
rect -192 -3548 -152 48
rect -140 15 3432 36
rect -140 -3254 -119 15
rect -140 -3515 -119 -3396
rect 3411 -104 3432 15
rect 3411 -3515 3432 -246
rect -140 -3536 3432 -3515
rect 3444 -3548 3484 48
rect -192 -3588 3150 -3548
rect 3292 -3588 3484 -3548
use pad  pad_4
array 0 8 350 0 0 102
timestamp 1763591700
transform 0 -1 -129 1 0 -3131
box 85 -25 227 77
use pad  pad_5
array 0 8 350 0 0 102
timestamp 1763591700
transform 1 0 265 0 1 25
box 85 -25 227 77
use pad  pad_6
array 0 8 350 0 0 102
timestamp 1763591700
transform 0 1 3421 -1 0 -369
box 85 -25 227 77
use pad  pad_7
array 0 8 350 0 0 102
timestamp 1763591700
transform -1 0 3027 0 -1 -3525
box 85 -25 227 77
<< labels >>
rlabel metal1 -1 0 141 102 1 Vdd
rlabel metal1 3396 -246 3498 -104 3 GND
rlabel metal1 3150 -3602 3292 -3500 5 Vdd
rlabel metal1 -206 -3396 -104 -3254 7 GND
rlabel metal1 454 94 462 106 1 phi0
rlabel metal1 477 0 486 7 1 phi1
rlabel space 827 0 836 7 1 phi2
rlabel metal1 1154 94 1162 111 1 reset
rlabel space 1177 0 1186 7 1 reset
rlabel metal1 1504 94 1512 103 1 top_0
rlabel metal1 1854 96 1862 103 1 top_1
rlabel metal1 2204 96 2212 103 1 top_2
rlabel metal1 2554 96 2562 103 1 top_3
rlabel metal1 2904 96 2912 103 1 top_4
rlabel metal1 3254 96 3262 103 1 top_5
rlabel metal1 3487 -566 3499 -558 1 right_0
rlabel metal1 3487 -916 3499 -908 1 right_1
rlabel metal1 3487 -1266 3499 -1258 1 right_2
rlabel metal1 3487 -1616 3499 -1608 1 right_3
rlabel metal1 3487 -1966 3499 -1958 1 right_4
rlabel metal1 3487 -2316 3499 -2308 1 right_5
rlabel metal1 3487 -2666 3499 -2658 1 right_6
rlabel metal1 3487 -3016 3499 -3008 1 right_7
rlabel metal1 3487 -3366 3499 -3358 1 right_8
rlabel metal1 2830 -3603 2838 -3591 5 bottom_0
rlabel metal1 2480 -3603 2488 -3591 5 bottom_1
rlabel metal1 2130 -3603 2138 -3591 5 bottom_2
rlabel metal1 1780 -3603 1788 -3591 5 bottom_3
rlabel metal1 1430 -3603 1438 -3591 5 bottom_4
rlabel metal1 1080 -3603 1088 -3591 5 bottom_5
rlabel metal1 730 -3603 738 -3591 5 bottom_6
rlabel metal1 380 -3603 388 -3591 5 bottom_7
rlabel metal1 30 -3603 38 -3591 5 bottom_8
rlabel metal1 -207 -2942 -195 -2934 1 left_0
rlabel metal1 -207 -2592 -195 -2584 1 left_1
rlabel space -207 -2242 -195 -2234 1 left_2
rlabel metal1 -207 -1892 -195 -1884 1 left_3
rlabel metal1 -207 -1542 -195 -1534 1 left_4
rlabel metal1 -207 -1192 -195 -1184 1 left_5
rlabel metal1 -207 -842 -195 -834 1 left_6
rlabel metal1 -207 -492 -195 -484 1 left_7
rlabel metal1 -207 -142 -195 -134 1 left_8
rlabel metal1 1406 97 1414 103 1 top_0_oe
rlabel metal1 1756 97 1764 103 1 top_1_oe
rlabel metal1 2106 97 2114 103 1 top_2_oe
rlabel metal1 2456 97 2464 103 1 top_3_oe
rlabel metal1 2806 97 2814 103 1 top_4_oe
rlabel metal1 3156 97 3164 103 1 top_5_oe
rlabel metal1 3493 -468 3499 -460 1 right_0_oe
rlabel metal1 3493 -818 3499 -810 1 right_1_oe
rlabel metal1 3493 -1168 3499 -1160 1 right_2_oe
rlabel metal1 3493 -1518 3499 -1510 1 right_3_oe
rlabel metal1 3493 -1868 3499 -1860 1 right_4_oe
rlabel metal1 3493 -2218 3499 -2210 1 right_5_oe
rlabel metal1 3493 -2568 3499 -2560 1 right_6_oe
rlabel metal1 3493 -2918 3499 -2910 1 right_7_oe
rlabel metal1 3493 -3268 3499 -3260 1 right_8_oe
rlabel metal1 2928 -3603 2936 -3597 5 bottom_0_oe
rlabel metal1 2578 -3603 2586 -3597 5 bottom_1_oe
rlabel metal1 2228 -3603 2236 -3597 5 bottom_2_oe
rlabel metal1 1878 -3603 1886 -3597 5 bottom_3_oe
rlabel metal1 1528 -3603 1536 -3597 5 bottom_4_oe
rlabel metal1 1178 -3603 1186 -3597 5 bottom_5_oe
rlabel metal1 828 -3603 836 -3597 5 bottom_6_oe
rlabel metal1 478 -3603 486 -3597 5 bottom_7_oe
rlabel metal1 128 -3603 136 -3597 5 bottom_8_oe
rlabel metal1 -207 -3040 -201 -3032 1 left_0_oe
rlabel metal1 -207 -2690 -201 -2682 1 left_1_oe
rlabel metal1 -207 -2340 -201 -2332 1 left_2_oe
rlabel metal1 -207 -1990 -201 -1982 1 left_3_oe
rlabel metal1 -207 -1640 -201 -1632 1 left_4_oe
rlabel metal1 -207 -1290 -201 -1282 1 left_5_oe
rlabel metal1 -207 -940 -201 -932 1 left_6_oe
rlabel metal1 -207 -590 -201 -582 1 left_7_oe
rlabel metal1 -207 -240 -201 -232 1 left_8_oe
rlabel metal1 804 96 812 108 1 phi1
<< end >>
