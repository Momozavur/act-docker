magic
tech scmos
timestamp 1761284462
<< nwell >>
rect 54 -33 113 -5
<< pwell >>
rect 54 -57 113 -34
<< ntransistor >>
rect 66 -45 68 -40
rect 75 -45 77 -40
rect 93 -45 95 -40
rect 99 -45 101 -40
<< ptransistor >>
rect 66 -27 68 -17
rect 75 -27 77 -17
rect 93 -27 95 -17
rect 99 -27 101 -17
<< ndiffusion >>
rect 65 -45 66 -40
rect 68 -45 69 -40
rect 74 -45 75 -40
rect 77 -45 78 -40
rect 92 -45 93 -40
rect 95 -45 99 -40
rect 101 -45 102 -40
<< pdiffusion >>
rect 65 -27 66 -17
rect 68 -27 69 -17
rect 74 -27 75 -17
rect 77 -27 78 -17
rect 92 -27 93 -17
rect 95 -27 99 -17
rect 101 -27 102 -17
<< ndcontact >>
rect 60 -45 65 -40
rect 69 -45 74 -40
rect 78 -45 83 -40
rect 87 -45 92 -40
rect 102 -45 107 -40
<< pdcontact >>
rect 60 -27 65 -17
rect 78 -27 83 -17
rect 102 -27 107 -17
<< nsubstratendiff >>
rect 57 -13 62 -8
<< psubstratepcontact >>
rect 57 -54 69 -49
<< nsubstratencontact >>
rect 62 -13 75 -8
<< polysilicon >>
rect 54 -6 86 -5
rect 54 -7 91 -6
rect 54 -28 56 -7
rect 66 -17 68 -14
rect 75 -17 77 -14
rect 93 -17 95 -14
rect 99 -17 101 -14
rect 66 -28 68 -27
rect 54 -30 68 -28
rect 66 -40 68 -30
rect 75 -40 77 -27
rect 93 -31 95 -27
rect 99 -30 101 -27
rect 93 -40 95 -36
rect 99 -40 101 -37
rect 66 -48 68 -45
rect 75 -51 77 -45
rect 93 -48 95 -45
rect 99 -51 101 -45
rect 75 -53 101 -51
rect 78 -56 83 -53
<< polycontact >>
rect 86 -6 91 -1
rect 99 -14 104 -9
rect 78 -61 83 -56
<< metal1 >>
rect 91 -6 112 -1
rect 69 -17 74 -13
rect 78 -14 99 -9
rect 78 -17 83 -14
rect 107 -22 112 -6
rect 60 -31 65 -27
rect 60 -40 65 -36
rect 78 -40 83 -27
rect 102 -40 107 -27
rect 69 -49 74 -45
rect 87 -49 92 -45
rect 69 -52 92 -49
rect 74 -53 92 -52
<< m2contact >>
rect 60 -36 65 -31
<< pm12contact >>
rect 90 -36 95 -31
<< pdm12contact >>
rect 69 -27 74 -17
rect 87 -27 92 -17
<< metal2 >>
rect 74 -27 87 -17
rect 65 -36 90 -31
<< m123contact >>
rect 57 -13 62 -8
rect 69 -57 74 -52
rect 83 -61 88 -56
<< labels >>
rlabel polysilicon 67 -29 67 -29 1 in
rlabel metal1 105 -34 105 -34 1 out
rlabel polysilicon 76 -16 76 -16 1 c
rlabel nsubstratencontact 67 -11 67 -11 1 Vdd!
rlabel psubstratepcontact 67 -53 67 -53 1 GND!
<< end >>
