magic
tech scmos
timestamp 1761180946
<< nwell >>
rect 68 15 162 80
<< pwell >>
rect 68 -24 162 15
<< ntransistor >>
rect 85 -11 87 9
rect 95 -11 97 9
rect 105 -11 107 9
rect 116 -11 118 9
rect 144 -11 146 9
<< ptransistor >>
rect 85 24 87 64
rect 95 24 97 64
rect 105 24 107 64
rect 116 24 118 64
rect 144 24 146 64
<< ndiffusion >>
rect 79 -11 85 9
rect 87 -11 89 9
rect 94 -11 95 9
rect 97 -11 99 9
rect 104 -11 105 9
rect 107 -11 109 9
rect 114 -11 116 9
rect 118 -11 124 9
rect 140 -11 144 9
rect 146 -11 150 9
<< pdiffusion >>
rect 79 24 85 64
rect 87 24 95 64
rect 97 24 105 64
rect 107 24 116 64
rect 118 24 124 64
rect 140 24 144 64
rect 146 24 150 64
<< ndcontact >>
rect 74 -11 79 9
rect 89 -11 94 9
rect 99 -11 104 9
rect 109 -11 114 9
rect 124 -11 129 9
rect 135 -11 140 9
rect 150 -11 155 9
<< pdcontact >>
rect 74 24 79 64
rect 124 24 129 64
rect 135 24 140 64
rect 150 24 155 64
<< psubstratepcontact >>
rect 99 -21 104 -16
rect 135 -21 140 -16
<< nsubstratencontact >>
rect 99 69 104 74
rect 135 69 140 74
<< polysilicon >>
rect 85 64 87 67
rect 95 64 97 67
rect 105 64 107 67
rect 116 64 118 67
rect 144 64 146 67
rect 85 9 87 24
rect 95 9 97 24
rect 105 9 107 24
rect 116 9 118 24
rect 144 19 146 24
rect 144 9 146 14
rect 85 -14 87 -11
rect 95 -14 97 -11
rect 105 -14 107 -11
rect 116 -14 118 -11
rect 144 -14 146 -11
<< polycontact >>
rect 141 14 146 19
<< metal1 >>
rect 74 69 99 74
rect 104 69 135 74
rect 140 69 155 74
rect 74 64 79 69
rect 135 64 140 69
rect 124 19 129 24
rect 150 19 155 24
rect 89 14 141 19
rect 150 14 162 19
rect 89 9 94 14
rect 109 9 114 14
rect 150 9 155 14
rect 74 -16 79 -11
rect 99 -16 104 -11
rect 124 -16 129 -11
rect 135 -16 140 -11
rect 74 -21 99 -16
rect 104 -21 135 -16
rect 140 -21 155 -16
<< labels >>
rlabel nwell 85 64 88 67 1 a
rlabel nwell 95 64 98 67 1 b
rlabel nwell 105 64 108 67 1 c
rlabel nwell 115 64 118 67 1 d
rlabel metal1 150 69 155 74 1 Vdd!
rlabel metal1 150 -21 155 -16 1 GND!
rlabel metal1 157 14 162 19 7 out
<< end >>
