magic
tech scmos
timestamp 1761082932
<< nwell >>
rect 16 -34 75 -6
<< pwell >>
rect 16 -58 75 -35
<< ntransistor >>
rect 28 -46 30 -41
rect 37 -46 39 -41
rect 55 -46 57 -41
rect 61 -46 63 -41
<< ptransistor >>
rect 28 -28 30 -18
rect 37 -28 39 -18
rect 55 -28 57 -18
rect 61 -28 63 -18
<< ndiffusion >>
rect 27 -46 28 -41
rect 30 -46 31 -41
rect 36 -46 37 -41
rect 39 -46 40 -41
rect 54 -46 55 -41
rect 57 -46 61 -41
rect 63 -46 64 -41
<< pdiffusion >>
rect 27 -28 28 -18
rect 30 -28 31 -18
rect 36 -28 37 -18
rect 39 -28 40 -18
rect 54 -28 55 -18
rect 57 -28 61 -18
rect 63 -28 64 -18
<< ndcontact >>
rect 22 -46 27 -41
rect 31 -46 36 -41
rect 40 -46 45 -41
rect 49 -46 54 -41
rect 64 -46 69 -41
<< pdcontact >>
rect 22 -28 27 -18
rect 40 -28 45 -18
rect 64 -28 69 -18
<< nsubstratendiff >>
rect 19 -14 24 -9
<< psubstratepcontact >>
rect 19 -55 31 -50
<< nsubstratencontact >>
rect 24 -14 37 -9
<< polysilicon >>
rect 28 -18 30 -15
rect 37 -18 39 -15
rect 55 -18 57 -15
rect 61 -18 63 -15
rect 28 -29 30 -28
rect 16 -31 30 -29
rect 28 -41 30 -31
rect 37 -41 39 -28
rect 55 -32 57 -28
rect 61 -31 63 -28
rect 55 -41 57 -37
rect 61 -41 63 -38
rect 28 -49 30 -46
rect 37 -52 39 -46
rect 55 -49 57 -46
rect 61 -52 63 -46
rect 37 -54 63 -52
<< polycontact >>
rect 61 -15 66 -10
rect 63 -54 67 -49
<< metal1 >>
rect 31 -18 36 -14
rect 40 -15 61 -10
rect 40 -18 45 -15
rect 22 -32 27 -28
rect 22 -41 27 -37
rect 40 -41 45 -28
rect 64 -32 69 -28
rect 64 -37 75 -32
rect 64 -41 69 -37
rect 31 -50 36 -46
rect 49 -50 54 -46
rect 31 -53 54 -50
rect 36 -55 54 -53
rect 67 -53 72 -49
<< m2contact >>
rect 22 -37 27 -32
<< pm12contact >>
rect 52 -37 57 -32
<< pdm12contact >>
rect 31 -28 36 -18
rect 49 -28 54 -18
<< metal2 >>
rect 36 -28 49 -18
rect 27 -37 52 -32
<< m123contact >>
rect 19 -14 24 -9
rect 31 -58 36 -53
rect 67 -58 72 -53
<< labels >>
rlabel polysilicon 29 -30 29 -30 1 in
rlabel metal1 67 -35 67 -35 1 out
rlabel polysilicon 38 -17 38 -17 1 c
rlabel nsubstratencontact 29 -12 29 -12 1 Vdd!
rlabel psubstratepcontact 29 -54 29 -54 1 GND!
<< end >>
