magic
tech scmos
timestamp 1761015633
<< metal1 >>
rect -14 774 1 779
rect 75 712 76 717
rect 75 703 76 708
rect -14 668 1 673
rect 75 606 76 611
rect 75 597 76 602
rect -14 562 1 567
rect 75 500 76 505
rect 75 491 76 496
rect -14 456 1 461
rect 75 394 76 399
rect 75 385 76 390
rect -14 350 1 355
rect 75 288 76 293
rect 75 279 76 284
rect -14 244 1 249
rect 75 182 76 187
rect 75 173 76 178
rect -14 138 1 143
rect 75 76 76 81
rect 75 67 76 72
rect -14 32 1 37
rect 75 -30 76 -25
rect 75 -39 76 -34
<< metal2 >>
rect -14 -42 -9 806
<< metal3 >>
rect -3 -42 2 806
rect 6 -42 11 806
rect 24 -42 29 806
rect 70 -42 75 806
use reg_one  reg_one_0
timestamp 1761015633
transform 1 0 2 0 1 -17
box -11 -25 74 81
use reg_one  reg_one_1
timestamp 1761015633
transform 1 0 2 0 1 89
box -11 -25 74 81
use reg_one  reg_one_2
timestamp 1761015633
transform 1 0 2 0 1 195
box -11 -25 74 81
use reg_one  reg_one_3
timestamp 1761015633
transform 1 0 2 0 1 301
box -11 -25 74 81
use reg_one  reg_one_4
timestamp 1761015633
transform 1 0 2 0 1 407
box -11 -25 74 81
use reg_one  reg_one_5
timestamp 1761015633
transform 1 0 2 0 1 513
box -11 -25 74 81
use reg_one  reg_one_6
timestamp 1761015633
transform 1 0 2 0 1 619
box -11 -25 74 81
use reg_one  reg_one_7
timestamp 1761015633
transform 1 0 2 0 1 725
box -11 -25 74 81
<< labels >>
rlabel metal1 75 712 76 717 7 port00
rlabel metal1 75 703 76 708 7 port01
rlabel metal1 75 606 76 611 7 port10
rlabel metal1 75 597 76 602 7 port11
rlabel metal1 75 500 76 505 7 port20
rlabel metal1 75 491 76 496 7 port21
rlabel metal1 75 394 76 399 7 port30
rlabel metal1 75 385 76 390 7 port31
rlabel metal1 75 288 76 293 7 port40
rlabel metal1 75 279 76 284 7 port41
rlabel metal1 75 182 76 187 7 port50
rlabel metal1 75 173 76 178 7 port51
rlabel metal1 75 76 76 81 7 port60
rlabel metal1 75 67 76 72 7 port61
rlabel metal1 75 -30 76 -25 7 port70
rlabel metal1 75 -39 76 -34 7 port71
rlabel metal3 6 801 11 806 5 Vdd!
rlabel metal3 24 801 29 806 5 GND!
rlabel metal1 -2 774 1 779 3 in0
rlabel metal1 -2 668 1 673 3 in1
rlabel metal1 -2 562 1 567 3 in2
rlabel metal1 -2 456 1 461 3 in3
rlabel metal1 -2 350 1 355 3 in4
rlabel metal1 -2 244 1 249 3 in5
rlabel metal1 -2 138 1 143 3 in6
rlabel metal1 -2 32 1 37 3 in7
rlabel metal3 70 801 75 806 6 w
rlabel metal3 -3 801 2 806 5 r1
rlabel metal2 -14 801 -9 806 4 r0
<< end >>
