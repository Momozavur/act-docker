magic
tech scmos
timestamp 1765339832
<< pwell >>
rect -12 28 -7 33
rect 49 28 57 33
<< metal1 >>
rect -29 33 -24 37
rect 33 33 38 37
rect -112 2 -84 3
rect -107 -2 -84 2
rect -68 -5 -63 7
rect 1 0 7 5
rect 1 -13 6 0
rect -10 -26 7 -21
rect -10 -29 -7 -26
rect -112 -36 -84 -35
rect -107 -40 -84 -36
rect -60 -65 -55 -31
rect -29 -32 -7 -29
rect -29 -39 -24 -32
rect 56 -33 61 -11
rect -9 -38 2 -35
rect 22 -38 61 -33
rect -9 -41 -4 -38
rect -5 -65 4 -60
rect -107 -73 -24 -68
rect 22 -73 45 -68
<< m2contact >>
rect -109 25 -104 30
rect -89 28 -84 33
rect -68 28 -63 33
rect -7 28 -2 33
rect 55 28 60 33
rect -109 6 -104 11
rect 13 9 18 14
rect -52 0 -47 5
rect -9 -4 -4 1
rect -109 -13 -104 -8
rect -89 -10 -84 -5
rect -52 -26 -47 -21
rect -109 -32 -104 -27
rect -3 -35 2 -30
rect -49 -46 -44 -41
rect 42 -46 47 -41
rect -49 -65 -44 -60
rect 45 -73 50 -68
<< metal2 >>
rect -104 6 -98 11
rect -103 -8 -98 6
rect -84 5 -79 33
rect -63 28 -7 33
rect -2 28 55 33
rect -49 18 18 23
rect -49 14 -44 18
rect 13 14 18 18
rect -84 0 -52 5
rect -104 -13 -98 -8
rect -84 -21 -79 -5
rect -84 -26 -52 -21
rect -104 -32 -98 -27
rect -103 -59 -98 -32
rect -9 -30 -4 -4
rect 13 -16 18 9
rect 8 -21 18 -16
rect -9 -35 -3 -30
rect 8 -41 13 -21
rect -44 -46 42 -41
rect -103 -60 -83 -59
rect -103 -64 -49 -60
rect -88 -65 -49 -64
<< m123contact >>
rect -29 37 -24 42
rect 33 37 38 42
rect -112 -3 -107 2
rect -49 9 -44 14
rect -68 -10 -63 -5
rect -112 -41 -107 -36
rect -112 -73 -107 -68
use inv  inv_3
timestamp 1765001281
transform 0 1 11 -1 0 -48
box -10 -13 20 40
use inv  inv_2
timestamp 1765001281
transform 0 -1 -13 1 0 -58
box -10 -13 20 40
use inv  inv_0
timestamp 1765001281
transform 0 -1 -73 1 0 13
box -10 -13 20 40
use inv  inv_1
timestamp 1765001281
transform 0 -1 -73 1 0 -25
box -10 -13 20 40
use 2mux_nr  2mux_nr_0
timestamp 1765248526
transform 1 0 -28 0 1 6
box -32 -38 29 27
use 2mux_nr  2mux_nr_1
timestamp 1765248526
transform 1 0 34 0 1 6
box -32 -38 29 27
<< labels >>
rlabel metal2 -45 30 -45 30 1 GND!
rlabel m2contact 50 -73 50 -68 8 o
rlabel metal1 -29 37 -24 37 5 u
rlabel metal1 -112 -2 -112 3 3 au
rlabel metal1 -112 -41 -112 -35 3 ad
rlabel metal2 -85 -63 -85 -63 1 Vdd!
rlabel metal1 -112 -73 -112 -68 2 a
rlabel metal1 33 37 38 37 5 s
<< end >>
