magic
tech scmos
timestamp 1761084926
<< polysilicon >>
rect 0 391 2 393
rect 0 339 2 341
rect 0 287 2 289
rect 0 235 2 237
rect 0 183 2 185
rect 0 131 2 133
rect 0 79 2 81
rect 0 27 2 29
<< metal1 >>
rect 56 385 59 390
rect 56 333 59 338
rect 56 281 59 286
rect 56 229 59 234
rect 56 177 59 182
rect 56 125 59 130
rect 56 73 59 78
rect 56 21 59 26
<< metal3 >>
rect 3 0 8 416
rect 15 0 20 416
rect 51 0 56 416
use latch_one  latch_one_0
array 0 0 59 0 7 52
timestamp 1761082932
transform 1 0 -16 0 1 58
box 16 -58 75 -6
<< labels >>
rlabel polysilicon 0 339 2 341 3 in1
rlabel polysilicon 0 287 2 289 3 in2
rlabel polysilicon 0 235 2 237 3 in3
rlabel polysilicon 0 183 2 185 3 in4
rlabel polysilicon 0 79 2 81 3 in6
rlabel polysilicon 0 27 2 29 3 in7
rlabel polysilicon 0 131 2 133 3 in5
rlabel metal1 56 333 59 338 7 out1
rlabel metal1 56 281 59 286 7 out2
rlabel metal1 56 229 59 234 7 out3
rlabel metal1 56 177 59 182 7 out4
rlabel metal1 56 125 59 130 7 out5
rlabel metal1 56 73 59 78 7 out6
rlabel metal1 56 21 59 26 7 out7
rlabel metal3 15 413 20 416 5 GND!
rlabel metal3 3 413 8 416 5 Vdd!
rlabel metal3 51 413 56 416 5 c
rlabel polysilicon 0 391 2 393 3 in0
rlabel metal1 56 385 59 390 7 out0
<< end >>
