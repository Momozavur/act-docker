magic
tech scmos
timestamp 1765250278
<< metal1 >>
rect -90 738 -77 743
rect 76 738 79 743
rect -82 651 -77 738
rect -90 581 -77 586
rect 76 581 79 586
rect -82 495 -77 581
rect -90 424 -77 429
rect 76 424 79 429
rect -82 338 -77 424
rect -90 267 -77 272
rect 76 267 79 272
rect -82 181 -77 267
rect -90 110 -77 115
rect 76 110 79 115
rect -82 24 -77 110
rect -90 -47 -77 -42
rect 76 -47 79 -42
rect -82 -133 -77 -47
rect -90 -204 -77 -199
rect 76 -204 79 -199
rect -82 -290 -77 -204
rect -90 -361 -77 -356
rect 76 -361 79 -356
<< metal3 >>
rect -33 815 -28 853
rect -72 810 -28 815
rect -87 770 -77 775
rect -87 586 -82 770
rect -74 613 -62 618
rect -87 581 -77 586
rect -87 456 -77 461
rect -87 272 -82 456
rect -67 429 -62 613
rect -77 424 -62 429
rect -73 299 -62 304
rect -87 267 -77 272
rect -87 142 -77 147
rect -87 -42 -82 142
rect -67 115 -62 299
rect -73 110 -62 115
rect -73 -15 -62 -10
rect -87 -47 -77 -42
rect -87 -172 -77 -167
rect -87 -356 -82 -172
rect -67 -199 -62 -15
rect -73 -204 -62 -199
rect -33 -324 -28 810
rect -71 -329 -28 -324
rect -87 -361 -77 -356
rect -33 -361 -28 -329
rect -23 -361 -18 853
rect -3 -361 2 853
rect 48 -361 53 853
use shift_one  shift_one_7
timestamp 1765250278
transform 1 0 26 0 1 -288
box -113 -73 63 42
use shift_one  shift_one_6
timestamp 1765250278
transform 1 0 26 0 1 -131
box -113 -73 63 42
use shift_one  shift_one_5
timestamp 1765250278
transform 1 0 26 0 1 26
box -113 -73 63 42
use shift_one  shift_one_4
timestamp 1765250278
transform 1 0 26 0 1 183
box -113 -73 63 42
use shift_one  shift_one_2
timestamp 1765250278
transform 1 0 26 0 1 497
box -113 -73 63 42
use shift_one  shift_one_1
timestamp 1765250278
transform 1 0 26 0 1 654
box -113 -73 63 42
use shift_one  shift_one_0
timestamp 1765250278
transform 1 0 26 0 1 811
box -113 -73 63 42
use shift_one  shift_one_3
timestamp 1765250278
transform 1 0 26 0 1 340
box -113 -73 63 42
<< labels >>
rlabel metal3 -3 853 2 853 5 u
rlabel metal3 48 853 53 853 5 s
rlabel metal3 -21 823 -21 823 1 Vdd!
rlabel metal1 -90 738 -90 743 3 a0
rlabel metal1 77 738 79 743 7 o0
rlabel metal1 -90 581 -90 586 3 a1
rlabel metal1 77 581 79 586 7 o1
rlabel metal1 -90 424 -90 429 3 a2
rlabel metal1 77 424 79 429 7 o2
rlabel metal1 77 267 79 272 7 o3
rlabel metal1 -90 267 -90 272 3 a3
rlabel metal1 77 110 79 115 7 o4
rlabel metal1 -90 110 -90 115 3 a4
rlabel metal1 77 -47 79 -42 7 o5
rlabel metal1 -90 -47 -90 -42 3 a5
rlabel metal1 77 -204 79 -199 7 o6
rlabel metal1 -90 -204 -90 -199 3 a6
rlabel metal1 77 -361 79 -356 8 o7
rlabel metal1 -90 -361 -90 -356 2 a7
rlabel metal3 -31 842 -31 842 1 GND!
<< properties >>
string name shift_one_0
<< end >>
