magic
tech scmos
timestamp 1759377783
<< pwell >>
rect -2 0 1254 2
rect -2 -32 1246 0
<< polysilicon >>
rect -7 131 1225 133
rect -7 -35 -5 131
rect 99 123 101 131
rect 256 123 258 131
rect 413 123 415 131
rect 570 123 572 131
rect 727 123 729 131
rect 884 123 886 131
rect 1041 123 1043 131
rect 1198 123 1200 131
rect 110 121 126 123
rect 267 121 283 123
rect 424 121 440 123
rect 581 121 597 123
rect 738 121 754 123
rect 895 121 911 123
rect 1052 121 1068 123
rect 1209 121 1225 123
rect 53 65 65 67
rect 210 65 222 67
rect 367 65 379 67
rect 524 65 536 67
rect 681 65 693 67
rect 838 65 850 67
rect 995 65 1007 67
rect 1152 65 1164 67
rect 63 59 65 65
rect 220 59 222 65
rect 377 59 379 65
rect 534 59 536 65
rect 691 59 693 65
rect 848 59 850 65
rect 1005 59 1007 65
rect 1162 59 1164 65
rect 35 -35 37 -29
rect 150 -30 152 -6
rect 192 -30 194 -29
rect 150 -32 194 -30
rect 307 -30 309 -5
rect 349 -30 351 -29
rect 307 -32 351 -30
rect 464 -30 466 -6
rect 506 -30 508 -29
rect 464 -32 508 -30
rect 621 -30 623 -5
rect 663 -30 665 -29
rect 621 -32 665 -30
rect 778 -30 780 -6
rect 820 -30 822 -29
rect 778 -32 822 -30
rect 935 -30 937 -5
rect 977 -30 979 -29
rect 935 -32 979 -30
rect 1092 -30 1094 -6
rect 1134 -30 1136 -29
rect 1092 -32 1136 -30
rect -7 -37 37 -35
<< polycontact >>
rect 147 -6 152 -1
rect 304 -5 309 0
rect 461 -6 466 -1
rect 618 -5 623 0
rect 775 -6 780 -1
rect 932 -5 937 0
rect 1089 -6 1094 -1
<< metal1 >>
rect -7 125 63 130
rect 112 125 220 130
rect 269 125 377 130
rect 426 125 534 130
rect 583 125 691 130
rect 740 125 848 130
rect 897 125 1005 130
rect 1054 125 1162 130
rect -7 -32 -2 125
rect 14 62 19 67
rect 102 62 107 65
rect 259 62 264 65
rect 416 62 421 65
rect 573 62 578 65
rect 730 62 735 65
rect 887 62 892 65
rect 1044 62 1049 65
rect 1201 62 1206 65
rect 14 57 1206 62
rect 14 54 19 57
rect 171 54 176 57
rect 328 54 333 57
rect 485 54 490 57
rect 642 54 647 57
rect 799 54 804 57
rect 956 54 961 57
rect 1113 54 1118 57
rect 1248 -16 1259 -11
rect 24 -32 29 -29
rect 181 -32 186 -29
rect 338 -32 343 -29
rect 495 -32 500 -29
rect 652 -32 657 -29
rect 809 -32 814 -29
rect 966 -32 971 -29
rect 1123 -32 1128 -29
rect -7 -37 1128 -32
rect 1123 -40 1128 -37
<< m2contact >>
rect 72 85 77 90
rect 229 85 234 90
rect 386 85 391 90
rect 543 85 548 90
rect 700 85 705 90
rect 857 85 862 90
rect 1014 85 1019 90
rect 1171 85 1176 90
rect 124 -6 129 -1
rect 281 -6 286 -1
rect 438 -6 443 -1
rect 595 -6 600 -1
rect 752 -6 757 -1
rect 909 -6 914 -1
rect 1066 -6 1071 -1
rect 1223 -6 1228 -1
<< metal2 >>
rect 72 59 77 85
rect 229 58 234 85
rect 386 59 391 85
rect 543 59 548 85
rect 700 59 705 85
rect 857 59 862 85
rect 1014 59 1019 85
rect 1171 59 1176 85
rect 124 -40 129 -6
rect 281 -40 286 -6
rect 438 -40 443 -6
rect 595 -40 600 -6
rect 752 -40 757 -6
rect 909 -40 914 -6
rect 1066 -40 1071 -6
rect 1223 -35 1228 -6
use addsub_one  addsub_one_0
timestamp 1759363553
transform 1 0 -7 0 1 25
box 5 -57 162 37
use xor  xor_0
timestamp 1759371655
transform -1 0 178 0 -1 79
box 55 -54 122 17
use addsub_one  addsub_one_1
timestamp 1759363553
transform 1 0 150 0 1 25
box 5 -57 162 37
use xor  xor_1
timestamp 1759371655
transform -1 0 335 0 -1 79
box 55 -54 122 17
use addsub_one  addsub_one_2
timestamp 1759363553
transform 1 0 307 0 1 25
box 5 -57 162 37
use xor  xor_2
timestamp 1759371655
transform -1 0 492 0 -1 79
box 55 -54 122 17
use addsub_one  addsub_one_3
timestamp 1759363553
transform 1 0 464 0 1 25
box 5 -57 162 37
use xor  xor_3
timestamp 1759371655
transform -1 0 649 0 -1 79
box 55 -54 122 17
use addsub_one  addsub_one_4
timestamp 1759363553
transform 1 0 621 0 1 25
box 5 -57 162 37
use xor  xor_4
timestamp 1759371655
transform -1 0 806 0 -1 79
box 55 -54 122 17
use addsub_one  addsub_one_5
timestamp 1759363553
transform 1 0 778 0 1 25
box 5 -57 162 37
use xor  xor_5
timestamp 1759371655
transform -1 0 963 0 -1 79
box 55 -54 122 17
use addsub_one  addsub_one_6
timestamp 1759363553
transform 1 0 935 0 1 25
box 5 -57 162 37
use xor  xor_6
timestamp 1759371655
transform -1 0 1120 0 -1 79
box 55 -54 122 17
use addsub_one  addsub_one_7
timestamp 1759363553
transform 1 0 1092 0 1 25
box 5 -57 162 37
use xor  xor_7
timestamp 1759371655
transform -1 0 1277 0 -1 79
box 55 -54 122 17
<< labels >>
rlabel metal1 1254 -16 1259 -11 7 cout
rlabel metal2 124 -40 129 -37 1 s0
rlabel metal2 281 -40 286 -37 1 s1
rlabel metal2 438 -40 443 -37 1 s2
rlabel metal2 595 -40 600 -37 1 s3
rlabel metal2 752 -40 757 -37 1 s4
rlabel metal2 909 -40 914 -37 1 s5
rlabel metal2 1066 -40 1071 -37 1 s6
rlabel metal2 1223 -35 1228 -32 1 s7
rlabel metal1 14 62 19 67 5 Vdd!
rlabel polysilicon 1222 131 1225 133 5 cin
rlabel metal1 1123 -40 1128 -37 1 GND!
rlabel polysilicon 53 65 56 67 1 a0
rlabel polysilicon 1222 121 1225 123 1 b7
rlabel polysilicon 123 121 126 123 1 b0
rlabel polysilicon 210 65 213 67 1 a1
rlabel polysilicon 367 65 370 67 1 a2
rlabel polysilicon 524 65 527 67 1 a3
rlabel polysilicon 681 65 684 67 1 a4
rlabel polysilicon 838 65 841 67 1 a5
rlabel polysilicon 995 65 998 67 1 a6
rlabel polysilicon 1152 65 1155 67 1 a7
rlabel polysilicon 1065 121 1068 123 1 b6
rlabel polysilicon 908 121 911 123 1 b5
rlabel polysilicon 751 121 754 123 1 b4
rlabel polysilicon 594 121 597 123 1 b3
rlabel polysilicon 437 121 440 123 1 b2
rlabel polysilicon 280 121 283 123 1 b1
<< end >>
