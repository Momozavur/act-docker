magic
tech scmos
timestamp 1765000963
<< error_p >>
rect -32 1 -27 13
rect -20 1 -15 6
rect -13 3 -9 7
rect -20 0 -14 1
rect -14 -6 -9 -1
<< nwell >>
rect -27 1 1 27
rect -27 0 -20 1
rect -15 0 1 1
rect -27 -38 1 0
<< pwell >>
rect 1 -38 29 27
<< ntransistor >>
rect 8 11 15 13
rect 8 -11 15 -9
rect 8 -24 15 -22
<< ptransistor >>
rect -13 11 -6 13
rect -14 -11 -7 -9
rect -14 -24 -7 -22
<< ndiffusion >>
rect 8 13 15 16
rect 8 8 15 11
rect 8 -9 15 -6
rect 8 -14 15 -11
rect 8 -22 15 -19
rect 8 -27 15 -24
<< pdiffusion >>
rect -13 13 -6 16
rect -13 8 -6 11
rect -14 -9 -7 -6
rect -14 -14 -7 -11
rect -14 -22 -7 -19
rect -14 -27 -7 -24
<< ndcontact >>
rect 8 16 15 21
rect 8 3 15 8
rect 8 -6 15 -1
rect 8 -19 15 -14
rect 8 -32 15 -27
<< pdcontact >>
rect -13 16 -6 21
rect -13 3 -6 8
rect -14 -6 -7 -1
rect -14 -19 -7 -14
rect -14 -32 -7 -27
<< psubstratepcontact >>
rect 21 -5 26 22
<< nsubstratencontact >>
rect -24 8 -19 22
<< polysilicon >>
rect -17 11 -13 13
rect -6 11 -1 13
rect 4 11 8 13
rect 15 11 19 13
rect -17 3 -15 11
rect -22 1 -15 3
rect -22 -22 -20 1
rect 17 -9 19 11
rect -17 -11 -14 -9
rect -7 -11 -4 -9
rect 5 -11 8 -9
rect 15 -11 19 -9
rect -1 -15 1 -14
rect -1 -17 5 -15
rect 3 -22 5 -17
rect -22 -24 -14 -22
rect -7 -24 -4 -22
rect 3 -24 8 -22
rect 15 -24 18 -22
<< polycontact >>
rect -1 11 4 16
<< metal1 >>
rect -24 22 -19 27
rect -19 16 -13 21
rect -1 16 4 27
rect 21 22 26 27
rect 15 16 21 21
rect -24 3 -19 8
rect -6 3 -1 8
rect 4 3 8 8
rect -27 -6 -14 -1
rect -7 -6 8 -1
rect 21 -10 26 -5
rect -7 -19 8 -17
rect 15 -19 29 -14
rect -14 -22 15 -19
rect -27 -32 -14 -27
rect -7 -32 8 -27
<< m2contact >>
rect -1 3 4 8
<< pm12contact >>
rect -4 -14 1 -9
<< metal2 >>
rect -1 -9 4 3
rect 1 -14 4 -9
<< labels >>
rlabel metal1 -1 27 4 27 5 s
rlabel metal1 21 27 26 27 5 GND!
rlabel metal1 29 -19 29 -14 7 out
rlabel metal1 -24 27 -19 27 5 Vdd!
rlabel metal1 -27 -6 -27 -1 3 in1
rlabel metal1 -27 -32 -27 -27 3 in0
<< end >>
