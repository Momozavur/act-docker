magic
tech scmos
timestamp 1759282424
<< metal1 >>
rect -90 738 -77 743
rect 76 738 79 743
rect -82 690 -77 738
rect -90 620 -77 625
rect 76 620 79 625
rect -82 573 -77 620
rect -90 502 -77 507
rect 76 502 79 507
rect -82 455 -77 502
rect -90 384 -77 389
rect 76 384 79 389
rect -82 337 -77 384
rect -90 266 -77 271
rect 76 266 79 271
rect -82 219 -77 266
rect -90 148 -77 153
rect 76 148 79 153
rect -82 101 -77 148
rect -90 30 -77 35
rect 76 30 79 35
rect -82 -17 -77 30
rect -90 -88 -77 -83
rect 76 -88 79 -83
<< metal3 >>
rect -34 813 -29 853
rect -73 808 -29 813
rect -87 770 -77 775
rect -87 625 -82 770
rect -74 652 -62 657
rect -87 620 -77 625
rect -87 534 -77 539
rect -87 389 -82 534
rect -67 507 -62 652
rect -77 502 -62 507
rect -73 416 -62 421
rect -87 384 -77 389
rect -87 298 -77 303
rect -87 153 -82 298
rect -67 271 -62 416
rect -73 266 -62 271
rect -73 180 -62 185
rect -87 148 -77 153
rect -87 62 -77 67
rect -87 -83 -82 62
rect -67 35 -62 180
rect -73 30 -62 35
rect -34 -51 -29 808
rect -72 -56 -29 -51
rect -87 -88 -77 -83
rect -34 -88 -29 -56
rect -23 -88 -18 853
rect -3 -88 2 853
rect 48 -88 53 853
use ud_shift  ud_shift_7
timestamp 1759282424
transform 1 0 26 0 1 811
box -103 -73 50 42
use ud_shift  ud_shift_0
timestamp 1759282424
transform 1 0 26 0 1 -15
box -103 -73 50 42
use ud_shift  ud_shift_1
timestamp 1759282424
transform 1 0 26 0 1 103
box -103 -73 50 42
use ud_shift  ud_shift_2
timestamp 1759282424
transform 1 0 26 0 1 221
box -103 -73 50 42
use ud_shift  ud_shift_3
timestamp 1759282424
transform 1 0 26 0 1 339
box -103 -73 50 42
use ud_shift  ud_shift_4
timestamp 1759282424
transform 1 0 26 0 1 457
box -103 -73 50 42
use ud_shift  ud_shift_5
timestamp 1759282424
transform 1 0 26 0 1 575
box -103 -73 50 42
use ud_shift  ud_shift_6
timestamp 1759282424
transform 1 0 26 0 1 693
box -103 -73 50 42
<< labels >>
rlabel metal3 -3 853 2 853 5 u
rlabel metal3 48 853 53 853 5 s
rlabel metal3 -32 842 -32 842 1 GND!
rlabel metal3 -21 823 -21 823 1 Vdd!
rlabel metal1 -90 -88 -90 -83 2 a7
rlabel metal1 -90 30 -90 35 3 a6
rlabel metal1 -90 738 -90 743 3 a0
rlabel metal1 -90 620 -90 625 3 a1
rlabel metal1 -90 502 -90 507 3 a2
rlabel metal1 -90 384 -90 389 3 a3
rlabel metal1 -90 266 -90 271 3 a4
rlabel metal1 -90 148 -90 153 3 a5
rlabel metal1 77 738 79 743 7 o0
rlabel metal1 77 620 79 625 7 o1
rlabel metal1 77 502 79 507 7 o2
rlabel metal1 77 384 79 389 7 o3
rlabel metal1 77 266 79 271 7 o4
rlabel metal1 77 148 79 153 7 o5
rlabel metal1 77 30 79 35 7 o6
rlabel metal1 77 -88 79 -83 8 o7
<< end >>
