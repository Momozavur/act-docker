magic
tech scmos
timestamp 1765741251
<< polysilicon >>
rect 182 26 184 35
rect 193 26 195 35
rect 171 -35 173 -9
rect 182 -35 184 -26
rect 193 -35 195 -26
rect 171 -96 173 -70
rect 182 -96 184 -87
rect 193 -96 195 -87
rect 171 -157 173 -131
rect 182 -157 184 -148
rect 193 -157 195 -148
<< polycontact >>
rect 181 35 186 40
rect 181 -26 186 -21
rect 181 -87 186 -82
rect 181 -148 186 -143
rect 166 -180 171 -175
<< metal1 >>
rect 74 -73 79 -47
rect 114 -73 119 40
rect 74 -78 119 -73
rect 114 -82 119 -78
rect 74 -125 79 -115
rect 114 -143 119 -87
rect 124 -11 129 40
rect 124 -110 129 -16
rect 124 -143 129 -115
rect 134 -21 139 35
rect 134 -47 139 -26
rect 134 -138 139 -52
rect 144 35 181 40
rect 144 -82 149 35
rect 186 3 191 8
rect 154 -21 159 -16
rect 154 -26 181 -21
rect 186 -58 191 -53
rect 144 -87 181 -82
rect 144 -120 149 -87
rect 186 -119 191 -114
rect 144 -138 149 -125
rect 124 -148 181 -143
rect 156 -180 166 -175
rect 186 -180 191 -175
<< m2contact >>
rect 104 -28 109 -23
rect 104 -52 109 -47
rect 104 -70 109 -65
rect 114 -87 119 -82
rect 104 -101 109 -96
rect 74 -115 79 -110
rect 104 -125 109 -120
rect 104 -143 109 -138
rect 114 -148 119 -143
rect 124 -16 129 -11
rect 124 -115 129 -110
rect 134 35 139 40
rect 134 -26 139 -21
rect 134 -52 139 -47
rect 202 27 207 32
rect 154 -16 159 -11
rect 212 -15 217 -10
rect 159 -35 164 -30
rect 202 -34 207 -29
rect 159 -76 164 -71
rect 212 -76 217 -71
rect 159 -96 164 -91
rect 202 -95 207 -90
rect 144 -125 149 -120
rect 159 -137 164 -132
rect 212 -137 217 -132
rect 202 -156 207 -151
rect 212 -198 217 -193
<< pm12contact >>
rect 191 35 196 40
rect 191 -26 196 -21
rect 191 -87 196 -82
rect 191 -148 196 -143
<< metal2 >>
rect 139 35 191 40
rect 202 32 207 39
rect 129 -16 154 -11
rect 139 -26 191 -21
rect 104 -30 109 -28
rect 202 -29 207 27
rect 104 -35 159 -30
rect 109 -52 134 -47
rect 104 -71 109 -70
rect 104 -76 159 -71
rect 119 -87 191 -82
rect 202 -90 207 -34
rect 104 -96 159 -91
rect 79 -115 124 -110
rect 109 -125 144 -120
rect 104 -137 159 -132
rect 104 -138 109 -137
rect 119 -148 191 -143
rect 202 -151 207 -95
rect 202 -205 207 -156
rect 212 -10 217 39
rect 212 -71 217 -15
rect 212 -132 217 -76
rect 212 -193 217 -137
rect 212 -205 217 -198
use 3nand  3nand_3
timestamp 1765694390
transform 1 0 86 0 1 -231
box 72 30 122 83
use 3nand  3nand_2
timestamp 1765694390
transform 1 0 86 0 1 -170
box 72 30 122 83
use inv2  inv2_1
timestamp 1765338958
transform 1 0 89 0 1 -133
box -10 -13 20 40
use decoder_nor2  decoder_nor2_2
timestamp 1765740216
transform 1 0 133 0 1 -229
box 68 24 149 85
use decoder_nor2  decoder_nor2_3
timestamp 1765740216
transform 1 0 133 0 1 -168
box 68 24 149 85
use 3nand  3nand_1
timestamp 1765694390
transform 1 0 86 0 1 -109
box 72 30 122 83
use inv2  inv2_0
timestamp 1765338958
transform 1 0 89 0 1 -60
box -10 -13 20 40
use decoder_nor2  decoder_nor2_1
timestamp 1765740216
transform 1 0 133 0 1 -107
box 68 24 149 85
use 3nand  3nand_0
timestamp 1765694390
transform 1 0 86 0 1 -48
box 72 30 122 83
use decoder_nor2  decoder_nor2_0
timestamp 1765740216
transform 1 0 133 0 1 -46
box 68 24 149 85
<< labels >>
rlabel metal2 202 35 207 39 5 Vdd!
rlabel metal2 212 35 217 39 5 GND!
rlabel metal1 186 3 191 8 1 out1
rlabel metal1 186 -58 191 -53 1 out2
rlabel metal1 186 -119 191 -114 1 out3
rlabel metal1 186 -180 191 -175 1 out4
rlabel metal1 74 -52 79 -47 3 in1
rlabel metal1 74 -125 79 -120 3 in2
rlabel metal1 156 -180 161 -175 1 e
<< end >>
