magic
tech scmos
timestamp 1765773944
<< pwell >>
rect 1489 1638 1494 1643
rect 1234 1616 1235 1625
<< polysilicon >>
rect 1298 1802 1300 1815
rect 1309 1802 1311 1815
<< polycontact >>
rect 1832 1790 1837 1795
rect 2332 1790 2337 1795
<< metal1 >>
rect 2644 3285 2649 3291
rect 2460 3134 2465 3139
rect 2470 3087 2475 3092
rect 2380 2595 2385 2600
rect 2360 2546 2365 2551
rect 2608 2257 2617 2266
rect 2608 2248 2660 2257
rect 1253 1758 1258 1784
rect 1805 1769 1814 1774
rect 2305 1769 2316 1774
rect 1253 1753 1278 1758
rect 1273 1634 1278 1753
rect 1286 1727 1291 1762
rect 1805 1729 1810 1769
rect 1805 1724 1816 1729
rect 1835 1725 1840 1732
rect 2305 1729 2310 1769
rect 2609 1737 2618 1764
rect 2305 1724 2316 1729
rect 2335 1722 2340 1737
rect 2609 1732 2640 1737
rect 2651 1732 2660 2248
rect 2611 1729 2616 1732
rect 2653 1728 2658 1732
rect 351 1561 356 1566
rect 3130 1535 3135 1540
rect 3254 1535 3259 1540
rect 351 1385 356 1390
rect 3130 1359 3135 1364
rect 3254 1359 3259 1364
rect 351 1209 356 1214
rect 3130 1183 3135 1188
rect 3254 1183 3259 1188
rect 351 1033 356 1038
rect 3130 1007 3135 1012
rect 3254 1007 3259 1012
rect 351 857 356 862
rect 3130 831 3135 836
rect 3254 831 3259 836
rect 351 681 356 686
rect 3130 655 3135 660
rect 3254 655 3259 660
rect 351 505 356 510
rect 3130 479 3135 484
rect 3254 479 3259 484
rect 351 329 356 334
rect 3130 303 3135 308
rect 3254 303 3259 308
<< m2contact >>
rect 2608 2266 2617 2275
rect 1317 1799 1322 1804
rect 2609 1764 2618 1773
rect 1853 1716 1858 1721
rect 1489 1638 1494 1643
rect 1959 1523 1964 1528
rect 1959 1347 1964 1352
rect 1959 1171 1964 1176
rect 1959 995 1964 1000
rect 1959 819 1964 824
rect 1959 643 1964 648
rect 1959 467 1964 472
rect 1959 291 1964 296
<< pm12contact >>
rect 1296 1815 1301 1820
rect 1309 1815 1314 1820
<< metal2 >>
rect 2598 2225 2603 2232
rect 1317 1754 1322 1799
rect 1848 1770 1862 1775
rect 2348 1770 2362 1775
rect 2594 1773 2603 2225
rect 1848 1716 1853 1770
rect 2348 1716 2353 1770
rect 2594 1764 2609 1773
rect 2681 1764 2690 2214
rect 2699 2205 2708 2222
rect 2699 1764 2708 2196
rect 2717 2187 2726 2222
rect 2717 1764 2726 2178
rect 2735 2169 2744 2222
rect 2735 1764 2744 2160
rect 2763 2151 2772 2222
rect 2763 1764 2772 2142
rect 2781 2133 2790 2222
rect 2781 1764 2790 2124
rect 2799 2115 2808 2222
rect 2799 1764 2808 2106
rect 2817 2097 2826 2222
rect 2817 1764 2826 2088
rect 2845 2079 2854 2222
rect 2845 1764 2854 2070
rect 2863 2061 2872 2222
rect 2863 1764 2872 2052
rect 2881 2043 2890 2222
rect 2881 1764 2890 2034
rect 2899 2025 2908 2222
rect 2899 1764 2908 2016
rect 2927 2007 2936 2222
rect 2927 1764 2936 1998
rect 2945 1989 2954 2222
rect 2945 1764 2954 1980
rect 2963 1971 2972 2222
rect 2963 1764 2972 1962
rect 2981 1953 2990 2222
rect 2981 1764 2990 1944
rect 3009 1935 3018 2222
rect 3009 1755 3018 1926
rect 3027 1917 3036 2222
rect 3027 1765 3036 1908
rect 3045 1899 3054 2222
rect 2384 1746 3018 1755
rect 3045 1737 3054 1890
rect 3063 1881 3072 2222
rect 3063 1764 3072 1872
rect 3091 1863 3100 2222
rect 3091 1764 3100 1854
rect 3109 1845 3118 2222
rect 3109 1764 3118 1836
rect 3127 1827 3136 2222
rect 3127 1764 3136 1818
rect 3145 1809 3154 2222
rect 3145 1764 3154 1800
rect 3173 1791 3182 2222
rect 3173 1764 3182 1782
rect 3189 1773 3198 2222
rect 3209 1764 3218 2222
rect 3227 1764 3236 2222
rect 3000 1728 3054 1737
rect 3000 1697 3009 1728
rect 2364 1688 3009 1697
rect 715 1612 782 1617
rect 1452 1612 1457 1616
rect 1559 1612 1564 1616
rect 1666 1612 1671 1616
rect 2364 1617 2373 1688
rect 1866 1612 1871 1615
rect 2366 1615 2373 1617
rect 2366 1612 2371 1615
rect 2473 1612 2478 1616
rect 2666 1612 2671 1616
rect 804 1611 864 1612
rect 804 1607 859 1611
rect 2661 1607 2671 1612
rect 3000 1608 3009 1688
<< m3contact >>
rect 2681 2214 2690 2223
rect 2699 2196 2708 2205
rect 2717 2178 2726 2187
rect 2735 2160 2744 2169
rect 2763 2142 2772 2151
rect 2781 2124 2790 2133
rect 2799 2106 2808 2115
rect 2817 2088 2826 2097
rect 2845 2070 2854 2079
rect 2863 2052 2872 2061
rect 2881 2034 2890 2043
rect 2899 2016 2908 2025
rect 2927 1998 2936 2007
rect 2945 1980 2954 1989
rect 2963 1962 2972 1971
rect 2981 1944 2990 1953
rect 3009 1926 3018 1935
rect 3027 1908 3036 1917
rect 3045 1890 3054 1899
rect 2375 1746 2384 1755
rect 3063 1872 3072 1881
rect 3091 1854 3100 1863
rect 3109 1836 3118 1845
rect 3127 1818 3136 1827
rect 3145 1800 3154 1809
rect 3173 1782 3182 1791
rect 3189 1764 3198 1773
rect 1559 1616 1564 1621
rect 1666 1616 1671 1621
<< m123contact >>
rect 2591 3285 2596 3291
rect 1832 1795 1837 1800
rect 2332 1795 2337 1800
rect 3002 1603 3007 1608
rect 1083 1563 1092 1572
<< metal3 >>
rect 2596 3285 2600 3291
rect 2591 2242 2600 3285
rect 1863 2232 2352 2242
rect 2363 2232 2600 2242
rect 411 2196 2699 2205
rect 411 1601 420 2196
rect 532 2178 2717 2187
rect 532 1576 541 2178
rect 885 2160 2735 2169
rect 885 1684 894 2160
rect 917 2142 2763 2151
rect 917 1684 926 2142
rect 951 2124 2781 2133
rect 951 1684 960 2124
rect 1057 2106 2799 2115
rect 1057 1706 1066 2106
rect 1083 2088 2817 2097
rect 986 1684 991 1689
rect 986 1653 991 1662
rect 715 1621 720 1626
rect 777 1621 782 1626
rect 936 1574 941 1653
rect 1083 1572 1092 2088
rect 1205 2070 2845 2079
rect 1205 1815 1214 2070
rect 1205 1634 1214 1810
rect 1225 2052 2863 2061
rect 1205 1625 1207 1634
rect 1225 1625 1234 2052
rect 1403 2034 2881 2043
rect 1403 1625 1412 2034
rect 1488 2016 2899 2025
rect 1488 1741 1497 2016
rect 1512 1998 2927 2007
rect 1512 1625 1521 1998
rect 1356 1616 1388 1621
rect 1403 1616 1436 1625
rect 1461 1616 1521 1625
rect 1534 1980 2945 1989
rect 1534 1616 1543 1980
rect 1641 1962 2963 1971
rect 1564 1616 1602 1621
rect 1641 1616 1650 1962
rect 1671 1616 1709 1621
rect 1748 1616 1757 1962
rect 1830 1944 2981 1953
rect 1830 1800 1842 1944
rect 1875 1926 3009 1935
rect 1875 1620 1884 1926
rect 1948 1908 3027 1917
rect 1429 1612 1434 1616
rect 1463 1612 1468 1616
rect 1536 1612 1541 1616
rect 1570 1612 1575 1616
rect 1597 1612 1602 1616
rect 1643 1612 1648 1616
rect 1677 1612 1682 1616
rect 1704 1611 1709 1616
rect 1750 1612 1755 1616
rect 1877 1615 1882 1620
rect 1948 1615 1957 1908
rect 2200 1890 3045 1899
rect 2200 1622 2209 1890
rect 2330 1872 3063 1881
rect 2330 1800 2342 1872
rect 2448 1854 3091 1863
rect 1950 1612 1955 1615
rect 2375 1620 2384 1746
rect 2200 1608 2209 1613
rect 2377 1612 2382 1620
rect 2448 1615 2457 1854
rect 2482 1836 3109 1845
rect 2482 1616 2491 1836
rect 2555 1818 3127 1827
rect 2555 1616 2564 1818
rect 2675 1800 3145 1809
rect 2675 1616 2684 1800
rect 2748 1782 3173 1791
rect 2748 1616 2757 1782
rect 3124 1764 3189 1773
rect 3198 1764 3258 1773
rect 2450 1612 2455 1615
rect 2484 1612 2489 1616
rect 2557 1612 2562 1616
rect 2677 1612 2682 1616
rect 2750 1612 2755 1616
rect 3124 1608 3133 1764
rect 3248 1608 3258 1764
rect 411 1568 416 1571
rect 536 1568 541 1571
rect 859 1561 864 1566
rect 1066 1561 1071 1566
rect 1327 1564 1332 1569
rect 2202 1568 2207 1574
rect 3002 1570 3007 1574
rect 3126 1571 3131 1575
rect 3250 1569 3255 1573
<< m234contact >>
rect 859 1606 864 1611
rect 878 1592 883 1597
rect 1296 1820 1301 1825
rect 1309 1810 1314 1815
rect 1465 1635 1470 1640
rect 1343 1616 1352 1625
rect 1866 1615 1871 1620
rect 1452 1605 1457 1610
rect 1490 1605 1495 1610
rect 2473 1607 2478 1612
rect 478 1546 483 1551
rect 878 1416 883 1421
rect 478 1370 483 1375
rect 878 1240 883 1245
rect 478 1194 483 1199
rect 878 1064 883 1069
rect 478 1018 483 1023
rect 878 888 883 893
rect 478 842 483 847
rect 878 712 883 717
rect 478 666 483 671
rect 878 536 883 541
rect 478 490 483 495
rect 878 360 883 365
rect 478 314 483 319
<< m4contact >>
rect 1852 2232 1863 2242
rect 2352 2232 2363 2242
rect 936 1653 941 1658
rect 981 1653 986 1658
rect 1205 1810 1214 1815
rect 1207 1625 1216 1634
rect 1225 1616 1234 1625
rect 1857 1738 1862 1743
rect 2357 1738 2362 1743
rect 2200 1613 2209 1622
rect 2511 1607 2516 1612
rect 469 1506 474 1511
rect 469 1330 474 1335
rect 469 1154 474 1159
rect 469 978 474 983
rect 469 802 474 807
rect 469 626 474 631
rect 469 450 474 455
rect 469 274 474 279
<< metal4 >>
rect 1301 1820 1470 1825
rect 1214 1810 1309 1815
rect 941 1653 981 1658
rect 1465 1640 1470 1820
rect 1852 1743 1863 2232
rect 2352 1743 2363 2232
rect 1852 1738 1857 1743
rect 1862 1738 1863 1743
rect 1234 1616 1343 1625
rect 1871 1613 2200 1622
rect 1457 1605 1490 1610
rect 2478 1607 2511 1612
use latch_one  latch_one_1
timestamp 1765002978
transform 0 -1 2296 -1 0 1779
box -11 -67 48 -12
use latch_one  latch_one_0
timestamp 1765002978
transform 0 -1 1796 -1 0 1779
box -11 -67 48 -12
use datapath  datapath_0
timestamp 1765751372
transform 1 0 431 0 1 -264
box -81 532 2885 2021
use 2and  2and_0
timestamp 1765747547
transform -1 0 1396 0 1 1729
box 68 29 138 82
use rom  rom_0
timestamp 1765759847
transform 1 0 2676 0 1 3129
box -350 -907 584 162
use ring  ring_0
timestamp 1765052771
transform 1 0 178 0 1 3594
box -207 -3603 3499 111
<< labels >>
rlabel metal1 351 1561 356 1566 3 data_out0
rlabel metal1 351 1385 356 1390 3 data_out1
rlabel metal1 351 1209 356 1214 3 data_out2
rlabel metal1 351 1033 356 1038 3 data_out3
rlabel metal1 351 857 356 862 3 data_out4
rlabel metal1 351 681 356 686 3 data_out5
rlabel metal1 351 505 356 510 3 data_out6
rlabel metal1 351 329 356 334 3 data_out7
rlabel m234contact 478 314 483 319 1 data_in7
rlabel m234contact 478 490 483 495 1 data_in6
rlabel m234contact 478 666 483 671 1 data_in5
rlabel m234contact 478 842 483 847 1 data_in4
rlabel m234contact 478 1018 483 1023 1 data_in3
rlabel m234contact 478 1194 483 1199 1 data_in2
rlabel m234contact 478 1370 483 1375 1 data_in1
rlabel m234contact 478 1546 483 1551 1 data_in0
rlabel metal2 3209 2045 3218 2054 1 r_-w
rlabel metal1 3254 1359 3259 1364 1 addr_out9
rlabel metal1 3254 1535 3259 1540 1 addr_out8
rlabel metal1 3254 1183 3259 1188 1 addr_out10
rlabel metal1 3254 1007 3259 1012 1 addr_out11
rlabel metal1 3254 831 3259 836 1 addr_out12
rlabel metal1 3254 655 3259 660 1 addr_out13
rlabel metal1 3254 479 3259 484 1 addr_out14
rlabel metal1 3254 303 3259 308 1 addr_out15
rlabel metal1 3130 1536 3135 1540 1 addr_out0
rlabel metal1 3130 1360 3135 1364 1 addr_out1
rlabel metal1 3130 1184 3135 1188 1 addr_out2
rlabel metal1 3130 1008 3135 1012 1 addr_out3
rlabel metal1 3130 832 3135 836 1 addr_out4
rlabel metal1 3130 656 3135 660 1 addr_out5
rlabel metal1 3130 480 3135 484 1 addr_out6
rlabel metal1 3130 304 3135 308 1 addr_out7
rlabel m3contact 2681 2214 2690 2223 1 IR_w
rlabel metal1 2360 2546 2365 2551 1 s3
rlabel metal1 2380 2595 2385 2600 1 s2
rlabel metal1 2460 3134 2465 3139 1 s1
rlabel metal1 2644 3285 2649 3291 1 phi1
rlabel metal1 2470 3087 2475 3092 1 s0
rlabel metal3 411 1568 416 1571 1 rd_dataout
rlabel metal3 536 1568 541 1571 1 ld_datain
rlabel metal3 715 1621 720 1626 1 os_u
rlabel metal3 777 1621 782 1626 1 os_s
rlabel metal3 859 1561 864 1566 1 ros
rlabel metal3 887 1684 892 1689 1 fb_g3
rlabel metal3 919 1684 924 1689 1 fb_g2
rlabel metal3 953 1684 958 1689 1 fb_g1
rlabel metal3 986 1684 991 1689 1 fb_g0
rlabel metal3 1066 1561 1071 1566 1 rfb
rlabel m123contact 1087 1565 1092 1570 1 as_sub
rlabel metal1 1273 1634 1278 1639 1 as_cin
rlabel m234contact 1345 1616 1350 1621 1 A_r0
rlabel metal3 1356 1616 1361 1621 1 A_r1
rlabel metal3 1327 1564 1332 1569 1 ras
rlabel m234contact 878 1592 883 1597 1 ry0
rlabel m234contact 878 1416 883 1421 1 ry1
rlabel m234contact 878 1240 883 1245 1 ry2
rlabel m234contact 878 1064 883 1069 1 ry3
rlabel m234contact 878 888 883 893 1 ry4
rlabel m234contact 878 712 883 717 1 ry5
rlabel m234contact 878 536 883 541 1 ry6
rlabel m234contact 878 360 883 365 1 ry7
rlabel m4contact 469 1506 474 1511 1 rx0
rlabel m4contact 469 1330 474 1335 1 rx1
rlabel m4contact 469 1154 474 1159 1 rx2
rlabel m4contact 469 978 474 983 1 rx3
rlabel m4contact 469 802 474 807 1 rx4
rlabel m4contact 469 626 474 631 1 rx5
rlabel m4contact 469 450 474 455 1 rx6
rlabel m4contact 469 274 474 279 1 rx7
rlabel m2contact 1959 1523 1964 1526 1 rx_PCL0
rlabel m2contact 1959 1347 1964 1350 1 rx_PCL1
rlabel m2contact 1959 1171 1964 1174 1 rx_PCL2
rlabel m2contact 1959 995 1964 998 1 rx_PCL3
rlabel m2contact 1959 819 1964 822 1 rx_PCL4
rlabel m2contact 1959 643 1964 646 1 rx_PCL5
rlabel m2contact 1959 467 1964 470 1 rx_PCL6
rlabel m2contact 1959 291 1964 294 1 rx_PCL7
rlabel metal3 1429 1612 1434 1616 1 A_w
rlabel metal2 1452 1612 1457 1616 1 DB_r0
rlabel metal3 1463 1612 1468 1616 1 DB_r1
rlabel metal3 1536 1612 1541 1616 1 DB_w
rlabel metal2 1559 1612 1564 1616 1 X_r0
rlabel metal3 1570 1612 1575 1616 1 X_r1
rlabel metal3 1643 1612 1648 1616 1 X_w
rlabel metal2 1666 1612 1671 1616 1 Y_r0
rlabel metal3 1677 1612 1682 1616 1 Y_r1
rlabel metal3 1750 1612 1755 1616 1 Y_w
rlabel metal3 1876 1622 1881 1627 1 PCL_r1
rlabel metal2 1866 1612 1871 1615 1 PCL_r0
rlabel metal3 1950 1612 1955 1615 1 PCL_w
rlabel metal3 2202 1571 2207 1574 1 rPCplus1L
rlabel metal2 2366 1612 2371 1615 1 PCH_r0
rlabel metal3 2377 1612 2382 1615 1 PCH_r1
rlabel metal3 2450 1612 2455 1615 1 PCH_w
rlabel metal2 2473 1612 2478 1616 1 ABL_r0
rlabel metal3 2484 1612 2489 1616 1 ABL_r1
rlabel metal3 2557 1612 2562 1616 1 ABL_w
rlabel metal1 2635 1732 2640 1736 1 ABH_w_sel
rlabel metal2 2666 1612 2671 1616 1 ABH_r0
rlabel metal3 2677 1612 2682 1616 1 ABH_r1
rlabel metal3 2750 1612 2755 1616 1 ABH_w
rlabel metal3 3002 1570 3007 1574 1 rPCplus1H
rlabel metal3 3126 1572 3131 1575 1 rd_addrL
rlabel metal3 3250 1570 3255 1573 1 rd_addrH
rlabel metal1 2335 1729 2339 1732 1 PCH_w_sel
rlabel metal1 1835 1725 1840 1732 1 PCL_w_sel
rlabel m123contact 2591 3285 2596 3291 1 phi0
rlabel metal3 1491 1741 1496 1746 1 Cflag_w
rlabel m2contact 1489 1638 1494 1643 1 Cflag
rlabel space 177 3682 319 3696 1 Vdd!
rlabel space 632 3688 640 3700 1 phi0
rlabel space 982 3690 990 3702 1 phi1
rlabel space 1332 3688 1340 3705 1 reset
rlabel space -29 3452 -17 3460 1 r-w_
rlabel space -29 3102 -17 3110 1 d0
rlabel space -29 2752 -17 2760 1 d1
rlabel space -29 2402 -17 2410 1 d2
rlabel space -29 2052 -17 2060 1 d3
rlabel space -29 1702 -17 1710 1 d4
rlabel space -29 1352 -18 1360 1 d5
rlabel space -29 1002 -17 1010 1 d6
rlabel space -29 652 -17 660 1 d7
rlabel space -28 198 -14 340 1 GND!
rlabel space 558 -9 566 3 1 a15
rlabel space 908 -9 916 3 1 a14
rlabel space 1258 -9 1266 3 1 a13
rlabel space 1608 -9 1616 3 1 a12
rlabel space 1958 -9 1966 3 1 a11
rlabel space 2308 -9 2316 3 1 a10
rlabel space 2658 -9 2666 3 1 a9
rlabel space 3008 -9 3016 3 1 a8
rlabel space 3328 -8 3470 6 1 Vdd!
rlabel space 3665 228 3677 236 1 a7
rlabel space 3665 578 3677 586 1 a6
rlabel space 3665 928 3677 936 1 a5
rlabel space 3665 1278 3677 1286 1 a4
rlabel space 3665 1628 3677 1636 1 a3
rlabel space 3665 1978 3677 1986 1 a2
rlabel space 3665 2328 3677 2336 1 a1
rlabel space 3665 2678 3677 2686 1 a0
rlabel space 3662 3348 3676 3490 1 GND!
<< end >>
