magic
tech scmos
timestamp 1765002088
<< nwell >>
rect 55 -19 122 17
<< pwell >>
rect 55 -55 122 -20
<< ntransistor >>
rect 67 -31 69 -26
rect 87 -31 89 -26
rect 67 -42 69 -37
rect 77 -42 79 -37
rect 98 -42 100 -37
rect 107 -42 109 -37
<< ptransistor >>
rect 67 -1 69 4
rect 77 -1 79 4
rect 98 -1 100 4
rect 107 -1 109 4
rect 67 -11 69 -6
rect 87 -11 89 -6
<< ndiffusion >>
rect 66 -31 67 -26
rect 69 -31 70 -26
rect 86 -31 87 -26
rect 89 -31 91 -26
rect 66 -42 67 -37
rect 69 -42 77 -37
rect 79 -42 91 -37
rect 96 -42 98 -37
rect 100 -42 107 -37
rect 109 -42 111 -37
<< pdiffusion >>
rect 66 -1 67 4
rect 69 -1 70 4
rect 75 -1 77 4
rect 79 -1 81 4
rect 96 -1 98 4
rect 100 -1 101 4
rect 106 -1 107 4
rect 109 -1 111 4
rect 66 -11 67 -6
rect 69 -11 70 -6
rect 86 -11 87 -6
rect 89 -11 91 -6
<< ndcontact >>
rect 70 -31 75 -26
rect 81 -31 86 -26
rect 91 -31 96 -26
rect 61 -42 66 -37
rect 91 -42 96 -37
rect 111 -42 116 -37
<< pdcontact >>
rect 70 -1 75 4
rect 91 -1 96 4
rect 101 -1 106 4
rect 111 -1 116 4
rect 70 -11 75 -6
rect 81 -11 86 -6
rect 91 -11 96 -6
<< psubstratepcontact >>
rect 91 -52 96 -47
<< nsubstratencontact >>
rect 70 9 75 14
<< polysilicon >>
rect 67 4 69 7
rect 77 4 79 7
rect 98 4 100 7
rect 107 4 109 7
rect 67 -6 69 -1
rect 67 -26 69 -11
rect 67 -37 69 -31
rect 77 -33 79 -1
rect 87 -6 89 -3
rect 87 -26 89 -11
rect 87 -33 89 -31
rect 77 -35 89 -33
rect 77 -37 79 -35
rect 98 -37 100 -1
rect 107 -37 109 -1
rect 67 -45 69 -42
rect 77 -45 79 -42
rect 98 -45 100 -42
rect 107 -45 109 -42
<< polycontact >>
rect 93 -21 98 -16
<< metal1 >>
rect 70 4 75 9
rect 81 4 116 9
rect 70 -6 75 -1
rect 75 -11 81 -6
rect 91 -16 96 -11
rect 91 -21 93 -16
rect 91 -26 96 -21
rect 75 -31 81 -26
rect 61 -47 66 -42
rect 76 -47 81 -31
rect 101 -37 106 -1
rect 96 -42 106 -37
rect 111 -47 116 -42
rect 61 -52 91 -47
rect 96 -52 116 -47
<< pm12contact >>
rect 109 -21 114 -16
<< pdm12contact >>
rect 61 -1 66 4
rect 81 -1 86 4
rect 61 -11 66 -6
<< ndm12contact >>
rect 61 -31 66 -26
<< metal2 >>
rect 66 -1 81 4
rect 61 -16 66 -11
rect 61 -21 109 -16
rect 61 -26 66 -21
<< labels >>
rlabel polysilicon 77 -15 79 -13 1 b
rlabel metal1 101 -31 106 -26 1 out
rlabel polysilicon 67 -15 69 -13 1 a
rlabel nsubstratencontact 70 9 75 14 5 Vdd!
rlabel psubstratepcontact 91 -52 96 -47 1 GND!
<< end >>
