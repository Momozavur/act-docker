magic
tech scmos
timestamp 1758867764
<< nwell >>
rect -24 -38 1 27
<< pwell >>
rect 2 -38 27 27
<< ntransistor >>
rect 8 11 15 13
rect 8 -11 15 -9
rect 8 -24 15 -22
<< ptransistor >>
rect -12 11 -5 13
rect -12 -11 -5 -9
rect -12 -24 -5 -22
<< ndiffusion >>
rect 8 13 15 16
rect 8 8 15 11
rect 8 -9 15 -6
rect 8 -14 15 -11
rect 8 -22 15 -19
rect 8 -27 15 -24
<< pdiffusion >>
rect -12 13 -5 16
rect -12 8 -5 11
rect -12 -9 -5 -6
rect -12 -14 -5 -11
rect -7 -19 -5 -14
rect -12 -22 -5 -19
rect -12 -27 -5 -24
<< ndcontact >>
rect 8 16 15 21
rect 8 3 15 8
rect 8 -6 15 -1
rect 8 -19 15 -14
rect 8 -32 15 -27
<< pdcontact >>
rect -12 16 -5 21
rect -12 3 -5 8
rect -12 -6 -5 -1
rect -12 -19 -7 -14
rect -12 -32 -5 -27
<< psubstratepcontact >>
rect 19 -5 24 22
<< nsubstratencontact >>
rect -21 8 -16 22
<< polysilicon >>
rect -15 11 -12 13
rect -5 11 -1 13
rect 4 11 8 13
rect 15 11 18 13
rect -15 -3 -13 11
rect -20 -5 -13 -3
rect -20 -22 -18 -5
rect 16 -9 18 11
rect -15 -11 -12 -9
rect -5 -11 -4 -9
rect 5 -11 8 -9
rect 15 -11 18 -9
rect -1 -15 1 -14
rect -1 -17 7 -15
rect 5 -22 7 -17
rect -20 -24 -12 -22
rect -5 -24 -2 -22
rect 5 -24 8 -22
rect 15 -24 18 -22
<< polycontact >>
rect -1 11 4 16
<< metal1 >>
rect -21 22 -16 27
rect -16 16 -12 21
rect -1 16 4 27
rect 19 22 24 27
rect 15 16 19 21
rect -21 3 -16 8
rect -5 3 -1 8
rect 4 3 8 8
rect -24 -6 -12 -1
rect -5 -6 8 -1
rect 19 -10 24 -5
rect -7 -19 8 -17
rect 15 -19 27 -14
rect -12 -22 13 -19
rect -24 -32 -12 -27
rect -5 -32 8 -27
<< m2contact >>
rect -1 3 4 8
<< pm12contact >>
rect -4 -14 1 -9
<< metal2 >>
rect -1 -9 4 3
rect 1 -14 4 -9
<< labels >>
rlabel metal1 -1 27 4 27 5 s
rlabel metal1 -24 -6 -24 -1 3 in1
rlabel metal1 -24 -32 -24 -27 3 in0
rlabel metal1 -21 27 -16 27 5 Vdd!
rlabel metal1 27 -19 27 -14 7 out
rlabel metal1 19 27 24 27 5 GND!
<< end >>
