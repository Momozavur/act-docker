magic
tech scmos
timestamp 1765002646
<< labels >>
rlabel metal1 105 -34 105 -34 1 out
rlabel polysilicon 76 -16 76 -16 1 c
rlabel polysilicon 67 -30 67 -30 1 in
rlabel nsubstratencontact 67 -10 67 -10 1 Vdd!
rlabel psubstratepcontact 67 -55 67 -55 1 GND!
<< end >>
