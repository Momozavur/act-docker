magic
tech scmos
timestamp 1759345730
<< metal1 >>
rect -6 96 0 101
rect -6 45 0 50
rect 92 45 121 50
rect -6 -57 0 -52
rect -6 -108 0 -103
rect 92 -108 121 -103
rect -6 -210 0 -205
rect -6 -261 0 -256
rect 92 -261 121 -256
rect -6 -363 0 -358
rect -6 -414 0 -409
rect 92 -414 121 -409
rect -6 -516 0 -511
rect -6 -567 0 -562
rect 92 -567 121 -562
rect -6 -669 0 -664
rect -6 -720 0 -715
rect 92 -720 121 -715
rect -6 -822 0 -817
rect -6 -873 0 -868
rect 92 -873 121 -868
rect -6 -975 0 -970
rect -6 -1026 0 -1021
rect 92 -1026 121 -1021
<< m3contact >>
rect 44 76 55 81
rect 44 -77 55 -72
rect 44 -230 55 -225
rect 44 -383 55 -378
rect 44 -536 55 -531
rect 44 -689 55 -684
rect 44 -842 55 -837
rect 44 -995 55 -990
<< m123contact >>
rect -6 147 5 152
rect 27 147 38 152
rect 61 147 72 152
rect 94 147 105 152
rect 109 65 120 70
rect -6 -6 5 -1
rect 27 -6 38 -1
rect 61 -6 72 -1
rect 94 -6 105 -1
rect 109 -88 120 -83
rect -6 -159 5 -154
rect 27 -159 38 -154
rect 61 -159 72 -154
rect 94 -159 105 -154
rect 109 -241 120 -236
rect -6 -312 5 -307
rect 27 -312 38 -307
rect 61 -312 72 -307
rect 94 -312 105 -307
rect 109 -394 120 -389
rect -6 -465 5 -460
rect 27 -465 38 -460
rect 61 -465 72 -460
rect 94 -465 105 -460
rect 109 -547 120 -542
rect -6 -618 5 -613
rect 27 -618 38 -613
rect 61 -618 72 -613
rect 94 -618 105 -613
rect 109 -700 120 -695
rect -6 -771 5 -766
rect 27 -771 38 -766
rect 61 -771 72 -766
rect 94 -771 105 -766
rect 109 -853 120 -848
rect -6 -924 5 -919
rect 27 -924 38 -919
rect 61 -924 72 -919
rect 94 -924 105 -919
rect 109 -1006 120 -1001
<< metal3 >>
rect -6 -1 5 147
rect -6 -154 5 -6
rect -6 -307 5 -159
rect -6 -460 5 -312
rect -6 -613 5 -465
rect -6 -766 5 -618
rect -6 -919 5 -771
rect 27 -1 38 147
rect 27 -154 38 -6
rect 27 -307 38 -159
rect 27 -460 38 -312
rect 27 -613 38 -465
rect 27 -766 38 -618
rect 27 -919 38 -771
rect 44 -72 55 76
rect 44 -225 55 -77
rect 44 -378 55 -230
rect 44 -531 55 -383
rect 44 -684 55 -536
rect 44 -837 55 -689
rect 44 -990 55 -842
rect 61 -1 72 147
rect 61 -154 72 -6
rect 61 -307 72 -159
rect 61 -460 72 -312
rect 61 -613 72 -465
rect 61 -766 72 -618
rect 61 -919 72 -771
rect 94 -1 105 147
rect 94 -154 105 -6
rect 94 -307 105 -159
rect 94 -460 105 -312
rect 94 -613 105 -465
rect 94 -766 105 -618
rect 94 -919 105 -771
rect 109 -83 120 65
rect 109 -236 120 -88
rect 109 -389 120 -241
rect 109 -542 120 -394
rect 109 -695 120 -547
rect 109 -848 120 -700
rect 109 -1001 120 -853
use fblock_one  fblock_one_0
timestamp 1759303105
transform 1 0 -1 0 1 90
box -5 -68 125 85
use fblock_one  fblock_one_1
timestamp 1759303105
transform 1 0 -1 0 1 -63
box -5 -68 125 85
use fblock_one  fblock_one_2
timestamp 1759303105
transform 1 0 -1 0 1 -216
box -5 -68 125 85
use fblock_one  fblock_one_3
timestamp 1759303105
transform 1 0 -1 0 1 -369
box -5 -68 125 85
use fblock_one  fblock_one_4
timestamp 1759303105
transform 1 0 -1 0 1 -522
box -5 -68 125 85
use fblock_one  fblock_one_5
timestamp 1759303105
transform 1 0 -1 0 1 -675
box -5 -68 125 85
use fblock_one  fblock_one_6
timestamp 1759303105
transform 1 0 -1 0 1 -828
box -5 -68 125 85
use fblock_one  fblock_one_7
timestamp 1759303105
transform 1 0 -1 0 1 -981
box -5 -68 125 85
<< labels >>
rlabel m123contact -2 149 -2 149 3 g3
rlabel m123contact 32 148 32 148 1 g2
rlabel m123contact 65 149 65 149 1 g1
rlabel m123contact 99 149 99 149 1 g0
rlabel m123contact 115 67 115 67 1 Vdd!
rlabel m3contact 50 78 50 78 1 GND!
rlabel metal1 -6 45 0 50 3 a0
rlabel metal1 -6 96 0 101 3 b0
rlabel metal1 -6 -57 0 -52 3 b1
rlabel metal1 -6 -108 0 -103 3 a1
rlabel metal1 -6 -210 0 -205 3 b2
rlabel metal1 -6 -261 0 -256 3 a2
rlabel metal1 -6 -363 0 -358 3 b3
rlabel metal1 -6 -414 0 -409 3 a3
rlabel metal1 -6 -516 0 -511 3 b4
rlabel metal1 -6 -567 0 -562 3 a4
rlabel metal1 -6 -669 0 -664 3 b5
rlabel metal1 -6 -720 0 -715 3 a5
rlabel metal1 -6 -822 0 -817 3 b6
rlabel metal1 -6 -873 0 -868 3 a6
rlabel metal1 -6 -975 0 -970 3 b7
rlabel metal1 -6 -1026 0 -1021 3 a7
rlabel metal1 92 45 121 50 1 f0
rlabel metal1 92 -108 121 -103 1 f1
rlabel metal1 92 -261 121 -256 1 f2
rlabel metal1 92 -414 121 -409 1 f3
rlabel metal1 92 -567 121 -562 1 f4
rlabel metal1 92 -720 121 -715 1 f5
rlabel metal1 92 -873 121 -868 1 f6
rlabel metal1 92 -1026 121 -1021 1 f7
<< end >>
