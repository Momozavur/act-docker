magic
tech scmos
timestamp 1765765914
<< metal5 >>
rect 10 28 14 40
rect 28 36 32 40
rect 24 32 32 36
rect 36 36 58 40
rect 20 28 28 32
rect 10 24 24 28
rect 10 10 14 24
rect 20 20 28 24
rect 24 16 32 20
rect 28 10 32 16
rect 36 14 40 36
rect 54 14 58 36
rect 36 10 58 14
rect 62 14 66 40
rect 84 36 102 40
rect 84 28 88 36
rect 84 24 100 28
rect 84 14 88 24
rect 106 18 110 40
rect 120 18 124 40
rect 106 14 124 18
rect 62 10 80 14
rect 84 10 102 14
rect 110 10 120 14
<< end >>
