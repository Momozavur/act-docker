magic
tech scmos
timestamp 1765002646
<< nwell >>
rect 53 -33 113 -1
<< pwell >>
rect 53 -61 113 -33
<< ntransistor >>
rect 66 -46 68 -41
rect 75 -46 77 -41
rect 93 -46 95 -41
rect 99 -46 101 -41
<< ptransistor >>
rect 66 -27 68 -17
rect 75 -27 77 -17
rect 93 -27 95 -17
rect 99 -27 101 -17
<< ndiffusion >>
rect 65 -46 66 -41
rect 68 -46 69 -41
rect 74 -46 75 -41
rect 77 -46 78 -41
rect 92 -46 93 -41
rect 95 -46 99 -41
rect 101 -46 102 -41
<< pdiffusion >>
rect 65 -27 66 -17
rect 68 -27 69 -17
rect 74 -27 75 -17
rect 77 -27 78 -17
rect 92 -27 93 -17
rect 95 -27 99 -17
rect 101 -27 102 -17
<< ndcontact >>
rect 60 -46 65 -41
rect 69 -46 74 -41
rect 78 -46 83 -41
rect 87 -46 92 -41
rect 102 -46 107 -41
<< pdcontact >>
rect 60 -27 65 -17
rect 78 -27 83 -17
rect 102 -27 107 -17
<< nsubstratendiff >>
rect 57 -12 62 -7
<< psubstratepcontact >>
rect 57 -56 69 -51
<< nsubstratencontact >>
rect 62 -12 75 -7
<< polysilicon >>
rect 53 -5 86 -3
rect 53 -29 55 -5
rect 66 -17 68 -14
rect 75 -17 77 -14
rect 93 -17 95 -14
rect 99 -17 101 -14
rect 66 -29 68 -27
rect 53 -31 68 -29
rect 66 -41 68 -31
rect 75 -41 77 -27
rect 93 -31 95 -27
rect 99 -30 101 -27
rect 93 -41 95 -36
rect 99 -41 101 -37
rect 66 -49 68 -46
rect 75 -52 77 -46
rect 93 -49 95 -46
rect 99 -52 101 -46
rect 75 -54 101 -52
rect 78 -58 83 -54
<< polycontact >>
rect 86 -6 91 -1
rect 99 -14 104 -9
rect 78 -63 83 -58
<< metal1 >>
rect 91 -6 112 -1
rect 69 -17 74 -12
rect 78 -14 99 -9
rect 78 -17 83 -14
rect 107 -22 112 -6
rect 60 -31 65 -27
rect 60 -41 65 -36
rect 78 -41 83 -27
rect 102 -41 107 -27
rect 69 -51 74 -46
rect 87 -51 92 -46
rect 69 -54 92 -51
rect 74 -55 92 -54
<< m2contact >>
rect 60 -36 65 -31
<< pm12contact >>
rect 90 -36 95 -31
<< pdm12contact >>
rect 69 -27 74 -17
rect 87 -27 92 -17
<< metal2 >>
rect 74 -27 87 -17
rect 65 -36 90 -31
<< m123contact >>
rect 57 -12 62 -7
rect 69 -59 74 -54
rect 83 -63 88 -58
<< labels >>
rlabel metal1 105 -34 105 -34 1 out
rlabel polysilicon 76 -16 76 -16 1 c
rlabel polysilicon 67 -30 67 -30 1 in
rlabel nsubstratencontact 67 -10 67 -10 1 Vdd!
rlabel psubstratepcontact 67 -55 67 -55 1 GND!
<< end >>
