magic
tech scmos
timestamp 1765248240
<< error_s >>
rect 27 175 30 176
rect 61 175 63 176
rect 94 175 97 176
rect 67 167 69 168
rect 33 132 35 135
rect 8 131 35 132
rect 8 130 33 131
rect 73 130 98 132
rect 2 127 33 130
rect 69 127 98 130
rect -6 124 124 127
rect -6 123 24 124
rect 27 123 57 124
rect 61 123 91 124
rect 94 123 124 124
rect -1 122 13 123
rect 65 122 78 123
rect 20 120 21 121
rect 85 120 86 121
rect 21 115 26 120
rect 65 116 67 119
rect 86 115 91 120
rect 14 109 18 113
rect 22 109 27 114
rect 79 109 83 113
rect 87 109 92 114
rect 0 79 2 84
rect 8 79 33 81
rect 65 79 67 84
rect -1 76 33 79
rect -6 73 59 76
rect 64 74 90 77
rect 62 73 92 74
rect -6 71 92 73
rect 100 71 105 73
rect -1 70 13 71
rect 70 70 84 71
rect 20 69 21 70
rect 21 64 26 69
rect 14 58 18 62
rect 22 58 27 63
rect 0 28 2 33
rect 62 21 65 22
rect 27 18 30 19
rect 61 18 63 19
rect 94 18 97 19
rect 67 10 69 11
rect 33 -25 35 -22
rect 8 -26 35 -25
rect 8 -27 33 -26
rect 73 -27 98 -25
rect 2 -30 33 -27
rect 69 -30 98 -27
rect -6 -33 124 -30
rect -6 -34 24 -33
rect 27 -34 57 -33
rect 61 -34 91 -33
rect 94 -34 124 -33
rect -1 -35 13 -34
rect 65 -35 78 -34
rect 20 -37 21 -36
rect 85 -37 86 -36
rect 21 -42 26 -37
rect 65 -41 67 -38
rect 86 -42 91 -37
rect 14 -48 18 -44
rect 22 -48 27 -43
rect 79 -48 83 -44
rect 87 -48 92 -43
rect 0 -78 2 -73
rect 8 -78 33 -76
rect 65 -78 67 -73
rect -1 -81 33 -78
rect -6 -84 59 -81
rect 64 -83 90 -80
rect 62 -84 92 -83
rect -6 -86 92 -84
rect 100 -86 105 -84
rect -1 -87 13 -86
rect 70 -87 84 -86
rect 20 -88 21 -87
rect 21 -93 26 -88
rect 14 -99 18 -95
rect 22 -99 27 -94
rect 0 -129 2 -124
rect 62 -136 65 -135
rect 27 -139 30 -138
rect 61 -139 63 -138
rect 94 -139 97 -138
rect 67 -147 69 -146
rect 33 -182 35 -179
rect 8 -183 35 -182
rect 8 -184 33 -183
rect 73 -184 98 -182
rect 2 -187 33 -184
rect 69 -187 98 -184
rect -6 -190 124 -187
rect -6 -191 24 -190
rect 27 -191 57 -190
rect 61 -191 91 -190
rect 94 -191 124 -190
rect -1 -192 13 -191
rect 65 -192 78 -191
rect 20 -194 21 -193
rect 85 -194 86 -193
rect 21 -199 26 -194
rect 65 -198 67 -195
rect 86 -199 91 -194
rect 14 -205 18 -201
rect 22 -205 27 -200
rect 79 -205 83 -201
rect 87 -205 92 -200
rect 0 -235 2 -230
rect 8 -235 33 -233
rect 65 -235 67 -230
rect -1 -238 33 -235
rect -6 -241 59 -238
rect 64 -240 90 -237
rect 62 -241 92 -240
rect -6 -243 92 -241
rect 100 -243 105 -241
rect -1 -244 13 -243
rect 70 -244 84 -243
rect 20 -245 21 -244
rect 21 -250 26 -245
rect 14 -256 18 -252
rect 22 -256 27 -251
rect 0 -286 2 -281
rect 62 -293 65 -292
rect 27 -296 30 -295
rect 61 -296 63 -295
rect 94 -296 97 -295
rect 67 -304 69 -303
rect 33 -339 35 -336
rect 8 -340 35 -339
rect 8 -341 33 -340
rect 73 -341 98 -339
rect 2 -344 33 -341
rect 69 -344 98 -341
rect -6 -347 124 -344
rect -6 -348 24 -347
rect 27 -348 57 -347
rect 61 -348 91 -347
rect 94 -348 124 -347
rect -1 -349 13 -348
rect 65 -349 78 -348
rect 20 -351 21 -350
rect 85 -351 86 -350
rect 21 -356 26 -351
rect 65 -355 67 -352
rect 86 -356 91 -351
rect 14 -362 18 -358
rect 22 -362 27 -357
rect 79 -362 83 -358
rect 87 -362 92 -357
rect 0 -392 2 -387
rect 8 -392 33 -390
rect 65 -392 67 -387
rect -1 -395 33 -392
rect -6 -398 59 -395
rect 64 -397 90 -394
rect 62 -398 92 -397
rect -6 -400 92 -398
rect 100 -400 105 -398
rect -1 -401 13 -400
rect 70 -401 84 -400
rect 20 -402 21 -401
rect 21 -407 26 -402
rect 14 -413 18 -409
rect 22 -413 27 -408
rect 0 -443 2 -438
rect 62 -450 65 -449
rect 27 -453 30 -452
rect 61 -453 63 -452
rect 94 -453 97 -452
rect 67 -461 69 -460
rect 33 -496 35 -493
rect 8 -497 35 -496
rect 8 -498 33 -497
rect 73 -498 98 -496
rect 2 -501 33 -498
rect 69 -501 98 -498
rect -6 -504 124 -501
rect -6 -505 24 -504
rect 27 -505 57 -504
rect 61 -505 91 -504
rect 94 -505 124 -504
rect -1 -506 13 -505
rect 65 -506 78 -505
rect 20 -508 21 -507
rect 85 -508 86 -507
rect 21 -513 26 -508
rect 65 -512 67 -509
rect 86 -513 91 -508
rect 14 -519 18 -515
rect 22 -519 27 -514
rect 79 -519 83 -515
rect 87 -519 92 -514
rect 0 -549 2 -544
rect 8 -549 33 -547
rect 65 -549 67 -544
rect -1 -552 33 -549
rect -6 -555 59 -552
rect 64 -554 90 -551
rect 62 -555 92 -554
rect -6 -557 92 -555
rect 100 -557 105 -555
rect -1 -558 13 -557
rect 70 -558 84 -557
rect 20 -559 21 -558
rect 21 -564 26 -559
rect 14 -570 18 -566
rect 22 -570 27 -565
rect 0 -600 2 -595
rect 62 -607 65 -606
rect 27 -610 30 -609
rect 61 -610 63 -609
rect 94 -610 97 -609
rect 67 -618 69 -617
rect 33 -653 35 -650
rect 8 -654 35 -653
rect 8 -655 33 -654
rect 73 -655 98 -653
rect 2 -658 33 -655
rect 69 -658 98 -655
rect -6 -661 124 -658
rect -6 -662 24 -661
rect 27 -662 57 -661
rect 61 -662 91 -661
rect 94 -662 124 -661
rect -1 -663 13 -662
rect 65 -663 78 -662
rect 20 -665 21 -664
rect 85 -665 86 -664
rect 21 -670 26 -665
rect 65 -669 67 -666
rect 86 -670 91 -665
rect 14 -676 18 -672
rect 22 -676 27 -671
rect 79 -676 83 -672
rect 87 -676 92 -671
rect 0 -706 2 -701
rect 8 -706 33 -704
rect 65 -706 67 -701
rect -1 -709 33 -706
rect -6 -712 59 -709
rect 64 -711 90 -708
rect 62 -712 92 -711
rect -6 -714 92 -712
rect 100 -714 105 -712
rect -1 -715 13 -714
rect 70 -715 84 -714
rect 20 -716 21 -715
rect 21 -721 26 -716
rect 14 -727 18 -723
rect 22 -727 27 -722
rect 0 -757 2 -752
rect 62 -764 65 -763
rect 27 -767 30 -766
rect 61 -767 63 -766
rect 94 -767 97 -766
rect 67 -775 69 -774
rect 33 -810 35 -807
rect 8 -811 35 -810
rect 8 -812 33 -811
rect 73 -812 98 -810
rect 2 -815 33 -812
rect 69 -815 98 -812
rect -6 -818 124 -815
rect -6 -819 24 -818
rect 27 -819 57 -818
rect 61 -819 91 -818
rect 94 -819 124 -818
rect -1 -820 13 -819
rect 65 -820 78 -819
rect 20 -822 21 -821
rect 85 -822 86 -821
rect 21 -827 26 -822
rect 65 -826 67 -823
rect 86 -827 91 -822
rect 14 -833 18 -829
rect 22 -833 27 -828
rect 79 -833 83 -829
rect 87 -833 92 -828
rect 0 -863 2 -858
rect 8 -863 33 -861
rect 65 -863 67 -858
rect -1 -866 33 -863
rect -6 -869 59 -866
rect 64 -868 90 -865
rect 62 -869 92 -868
rect -6 -871 92 -869
rect 100 -871 105 -869
rect -1 -872 13 -871
rect 70 -872 84 -871
rect 20 -873 21 -872
rect 21 -878 26 -873
rect 14 -884 18 -880
rect 22 -884 27 -879
rect 0 -914 2 -909
rect 62 -921 65 -920
rect 27 -924 30 -923
rect 61 -924 63 -923
rect 94 -924 97 -923
rect 67 -932 69 -931
rect 33 -967 35 -964
rect 8 -968 35 -967
rect 8 -969 33 -968
rect 73 -969 98 -967
rect 2 -972 33 -969
rect 69 -972 98 -969
rect -6 -975 124 -972
rect -6 -976 24 -975
rect 27 -976 57 -975
rect 61 -976 91 -975
rect 94 -976 124 -975
rect -1 -977 13 -976
rect 65 -977 78 -976
rect 20 -979 21 -978
rect 85 -979 86 -978
rect 21 -984 26 -979
rect 65 -983 67 -980
rect 86 -984 91 -979
rect 14 -990 18 -986
rect 22 -990 27 -985
rect 79 -990 83 -986
rect 87 -990 92 -985
rect 0 -1020 2 -1015
rect 8 -1020 33 -1018
rect 65 -1020 67 -1015
rect -1 -1023 33 -1020
rect -6 -1026 59 -1023
rect 64 -1025 90 -1022
rect 62 -1026 92 -1025
rect -6 -1028 92 -1026
rect 100 -1028 105 -1026
rect -1 -1029 13 -1028
rect 70 -1029 84 -1028
rect 20 -1030 21 -1029
rect 21 -1035 26 -1030
rect 14 -1041 18 -1037
rect 22 -1041 27 -1036
rect 0 -1071 2 -1066
rect 62 -1078 65 -1077
<< metal1 >>
rect -6 96 0 101
rect -6 45 0 50
rect 92 45 121 50
rect -6 -61 0 -56
rect -6 -112 0 -107
rect 92 -112 121 -107
rect -6 -218 0 -213
rect -6 -269 0 -264
rect 92 -269 121 -264
rect -6 -375 0 -370
rect -6 -426 0 -421
rect 92 -426 121 -421
rect -6 -532 0 -527
rect -6 -583 0 -578
rect 92 -583 121 -578
rect -6 -689 0 -684
rect -6 -740 0 -735
rect 92 -740 121 -735
rect -6 -846 0 -841
rect -6 -897 0 -892
rect 92 -897 121 -892
rect -6 -1003 0 -998
rect -6 -1054 0 -1049
rect 92 -1054 121 -1049
<< m3contact >>
rect 44 76 55 81
rect 44 -81 55 -76
rect 44 -238 55 -233
rect 44 -395 55 -390
rect 44 -552 55 -547
rect 44 -709 55 -704
rect 44 -866 55 -861
rect 44 -1023 55 -1018
<< m123contact >>
rect -6 147 5 152
rect 27 147 38 152
rect 61 147 72 152
rect 94 147 105 152
rect 109 65 120 70
rect -6 -10 5 -5
rect 27 -10 38 -5
rect 61 -10 72 -5
rect 94 -10 105 -5
rect 109 -92 120 -87
rect -6 -167 5 -162
rect 27 -167 38 -162
rect 61 -167 72 -162
rect 94 -167 105 -162
rect 109 -249 120 -244
rect -6 -324 5 -319
rect 27 -324 38 -319
rect 61 -324 72 -319
rect 94 -324 105 -319
rect 109 -406 120 -401
rect -6 -481 5 -476
rect 27 -481 38 -476
rect 61 -481 72 -476
rect 94 -481 105 -476
rect 109 -563 120 -558
rect -6 -638 5 -633
rect 27 -638 38 -633
rect 61 -638 72 -633
rect 94 -638 105 -633
rect 109 -720 120 -715
rect -6 -795 5 -790
rect 27 -795 38 -790
rect 61 -795 72 -790
rect 94 -795 105 -790
rect 109 -877 120 -872
rect -6 -952 5 -947
rect 27 -952 38 -947
rect 61 -952 72 -947
rect 94 -952 105 -947
rect 109 -1034 120 -1029
<< metal3 >>
rect -6 -5 5 147
rect -6 -162 5 -10
rect -6 -319 5 -167
rect -6 -476 5 -324
rect -6 -633 5 -481
rect -6 -790 5 -638
rect -6 -947 5 -795
rect 27 -5 38 147
rect 27 -162 38 -10
rect 27 -319 38 -167
rect 27 -476 38 -324
rect 27 -633 38 -481
rect 27 -790 38 -638
rect 27 -947 38 -795
rect 44 81 55 106
rect 44 -76 55 76
rect 44 -233 55 -81
rect 44 -390 55 -238
rect 44 -547 55 -395
rect 44 -704 55 -552
rect 44 -861 55 -709
rect 44 -1018 55 -866
rect 61 -5 72 147
rect 61 -162 72 -10
rect 61 -319 72 -167
rect 61 -476 72 -324
rect 61 -633 72 -481
rect 61 -790 72 -638
rect 61 -947 72 -795
rect 94 -5 105 147
rect 94 -162 105 -10
rect 94 -319 105 -167
rect 94 -476 105 -324
rect 94 -633 105 -481
rect 94 -790 105 -638
rect 94 -947 105 -795
rect 109 -87 120 65
rect 109 -244 120 -92
rect 109 -401 120 -249
rect 109 -558 120 -406
rect 109 -715 120 -563
rect 109 -872 120 -720
rect 109 -1029 120 -877
use fblock_one  fblock_one_1
timestamp 1765248240
transform 1 0 -1 0 1 -67
box -5 -70 125 86
use fblock_one  fblock_one_2
timestamp 1765248240
transform 1 0 -1 0 1 -224
box -5 -70 125 86
use fblock_one  fblock_one_3
timestamp 1765248240
transform 1 0 -1 0 1 -381
box -5 -70 125 86
use fblock_one  fblock_one_4
timestamp 1765248240
transform 1 0 -1 0 1 -538
box -5 -70 125 86
use fblock_one  fblock_one_5
timestamp 1765248240
transform 1 0 -1 0 1 -695
box -5 -70 125 86
use fblock_one  fblock_one_6
timestamp 1765248240
transform 1 0 -1 0 1 -852
box -5 -70 125 86
use fblock_one  fblock_one_7
timestamp 1765248240
transform 1 0 -1 0 1 -1009
box -5 -70 125 86
use fblock_one  fblock_one_0
timestamp 1765248240
transform 1 0 -1 0 1 90
box -5 -70 125 86
<< labels >>
rlabel m123contact -2 149 -2 149 3 g3
rlabel m123contact 32 148 32 148 1 g2
rlabel m123contact 65 149 65 149 1 g1
rlabel m123contact 99 149 99 149 1 g0
rlabel m123contact 115 67 115 67 1 Vdd!
rlabel m3contact 50 78 50 78 1 GND!
rlabel metal1 -6 45 0 50 3 a0
rlabel metal1 -6 96 0 101 3 b0
rlabel metal1 92 45 121 50 1 f0
rlabel metal1 -6 -61 0 -56 3 b1
rlabel metal1 -6 -112 0 -107 3 a1
rlabel metal1 92 -112 121 -107 1 f1
rlabel metal1 -6 -218 0 -213 3 b2
rlabel metal1 -6 -269 0 -264 3 a2
rlabel metal1 92 -269 121 -264 1 f2
rlabel metal1 -6 -375 0 -370 3 b3
rlabel metal1 -6 -426 0 -421 3 a3
rlabel metal1 92 -426 121 -421 1 f3
rlabel metal1 92 -583 121 -578 1 f4
rlabel metal1 -6 -583 0 -578 3 a4
rlabel metal1 -6 -532 0 -527 3 b4
rlabel metal1 92 -740 121 -735 1 f5
rlabel metal1 -6 -740 0 -735 3 a5
rlabel metal1 -6 -689 0 -684 3 b5
rlabel metal1 92 -897 121 -892 1 f6
rlabel metal1 -6 -897 0 -892 3 a6
rlabel metal1 -6 -846 0 -841 3 b6
rlabel metal1 92 -1054 121 -1049 1 f7
rlabel metal1 -6 -1054 0 -1049 3 a7
rlabel metal1 -6 -1003 0 -998 3 b7
<< end >>
