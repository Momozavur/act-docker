magic
tech scmos
timestamp 1761179007
<< nwell >>
rect 68 15 162 80
<< pwell >>
rect 68 -24 162 15
<< ntransistor >>
rect 85 -11 88 9
rect 95 -11 98 9
rect 105 -11 108 9
rect 115 -11 118 9
rect 143 -11 147 9
<< ptransistor >>
rect 85 24 88 64
rect 95 24 98 64
rect 105 24 108 64
rect 115 24 118 64
rect 143 24 147 64
<< ndiffusion >>
rect 79 -11 85 9
rect 88 -11 89 9
rect 94 -11 95 9
rect 98 -11 99 9
rect 104 -11 105 9
rect 108 -11 109 9
rect 114 -11 115 9
rect 118 -11 124 9
rect 140 -11 143 9
rect 147 -11 150 9
<< pdiffusion >>
rect 79 24 85 64
rect 88 24 95 64
rect 98 24 105 64
rect 108 24 115 64
rect 118 24 124 64
rect 140 24 143 64
rect 147 24 150 64
<< ndcontact >>
rect 74 -11 79 9
rect 89 -11 94 9
rect 99 -11 104 9
rect 109 -11 114 9
rect 124 -11 129 9
rect 135 -11 140 9
rect 150 -11 155 9
<< pdcontact >>
rect 74 24 79 64
rect 124 24 129 64
rect 135 24 140 64
rect 150 24 155 64
<< psubstratepcontact >>
rect 99 -21 104 -16
<< nsubstratencontact >>
rect 99 69 104 74
<< polysilicon >>
rect 85 64 88 67
rect 95 64 98 67
rect 105 64 108 67
rect 115 64 118 67
rect 143 64 147 67
rect 85 9 88 24
rect 95 9 98 24
rect 105 9 108 24
rect 115 9 118 24
rect 143 19 147 24
rect 143 9 147 14
rect 85 -14 88 -11
rect 95 -14 98 -11
rect 105 -14 108 -11
rect 115 -14 118 -11
rect 143 -14 147 -11
<< polycontact >>
rect 142 14 147 19
<< metal1 >>
rect 74 69 99 74
rect 104 69 155 74
rect 74 64 79 69
rect 135 64 140 69
rect 150 64 155 69
rect 124 19 129 24
rect 150 19 155 24
rect 89 14 115 19
rect 118 14 142 19
rect 150 14 162 19
rect 89 9 94 14
rect 109 9 114 14
rect 150 9 155 14
rect 74 -16 79 -11
rect 99 -16 104 -11
rect 124 -16 129 -11
rect 135 -16 140 -11
rect 150 -16 155 -11
rect 74 -21 99 -16
rect 104 -21 155 -16
<< labels >>
rlabel polysilicon 85 64 88 67 1 a
rlabel polysilicon 95 64 98 67 1 b
rlabel polysilicon 105 64 108 67 1 c
rlabel polysilicon 115 64 118 67 1 d
rlabel metal1 150 69 155 74 1 Vdd!
rlabel metal1 150 -21 155 -16 1 GND!
rlabel metal1 157 14 162 19 7 out
<< end >>
