magic
tech scmos
timestamp 1765694390
<< nwell >>
rect 72 54 122 83
<< pwell >>
rect 72 30 122 53
<< ntransistor >>
rect 85 42 87 47
rect 96 42 98 47
rect 107 42 109 47
<< ptransistor >>
rect 85 61 87 71
rect 96 61 98 71
rect 107 61 109 71
<< ndiffusion >>
rect 83 42 85 47
rect 87 42 96 47
rect 98 42 107 47
rect 109 42 111 47
<< pdiffusion >>
rect 83 61 85 71
rect 87 61 89 71
rect 94 61 96 71
rect 98 61 100 71
rect 105 61 107 71
rect 109 61 111 71
<< ndcontact >>
rect 78 42 83 47
rect 111 42 116 47
<< pdcontact >>
rect 78 61 83 71
rect 89 61 94 71
rect 100 61 105 71
rect 111 61 116 71
<< psubstratepcontact >>
rect 100 33 105 38
<< nsubstratencontact >>
rect 100 75 105 80
<< polysilicon >>
rect 85 71 87 74
rect 96 71 98 74
rect 107 71 109 74
rect 85 47 87 61
rect 96 47 98 61
rect 107 47 109 61
rect 85 39 87 42
rect 96 39 98 42
rect 107 39 109 42
<< metal1 >>
rect 78 75 100 80
rect 105 75 122 80
rect 78 71 83 75
rect 100 71 105 75
rect 89 56 94 61
rect 111 56 116 61
rect 89 51 122 56
rect 111 47 116 51
rect 78 38 83 42
rect 78 33 100 38
rect 105 33 122 38
<< labels >>
rlabel polysilicon 85 72 87 74 1 a
rlabel polysilicon 96 72 98 74 1 b
rlabel metal1 117 33 122 38 7 GND!
rlabel metal1 117 75 122 80 7 Vdd!
rlabel polysilicon 107 72 109 74 1 c
rlabel metal1 117 51 122 56 7 out
<< end >>
