magic
tech scmos
timestamp 1765425687
<< polysilicon >>
rect 424 1804 425 1806
rect 424 1628 425 1630
rect 424 1452 425 1454
rect 424 1276 425 1278
rect 424 1100 425 1102
rect 424 924 425 926
rect 424 748 425 750
rect 424 572 425 574
<< polycontact >>
rect 477 1874 482 1879
rect -20 1800 -15 1805
rect 109 1800 114 1805
rect 326 1795 331 1800
rect 841 1796 846 1801
rect 477 1698 482 1703
rect -20 1624 -15 1629
rect 109 1624 114 1629
rect 326 1619 331 1624
rect 841 1620 846 1625
rect -20 1448 -15 1453
rect 109 1448 114 1453
rect 326 1443 331 1448
rect 841 1444 846 1449
rect -20 1272 -15 1277
rect 109 1272 114 1277
rect 326 1267 331 1272
rect 841 1268 846 1273
rect -20 1096 -15 1101
rect 109 1096 114 1101
rect 326 1091 331 1096
rect 841 1092 846 1097
rect -20 920 -15 925
rect 109 920 114 925
rect 326 915 331 920
rect 841 916 846 921
rect -20 744 -15 749
rect 109 744 114 749
rect 326 739 331 744
rect 841 740 846 745
rect -20 568 -15 573
rect 109 568 114 573
rect 326 563 331 568
rect 841 564 846 569
<< metal1 >>
rect -76 1825 -71 1830
rect 165 1825 170 1830
rect 309 1795 326 1800
rect 837 1796 841 1801
rect 837 1775 842 1796
rect 831 1770 842 1775
rect -76 1649 -71 1654
rect 165 1649 170 1654
rect 309 1619 326 1624
rect 837 1620 841 1625
rect 837 1599 842 1620
rect 831 1594 842 1599
rect -76 1473 -71 1478
rect 165 1473 170 1478
rect 309 1443 326 1448
rect 837 1444 841 1449
rect 837 1423 842 1444
rect 831 1418 842 1423
rect -76 1297 -71 1302
rect 165 1297 170 1302
rect 309 1267 326 1272
rect 837 1268 841 1273
rect 837 1247 842 1268
rect 831 1242 842 1247
rect -76 1121 -71 1126
rect 165 1121 170 1126
rect 309 1091 326 1096
rect 837 1092 841 1097
rect 837 1071 842 1092
rect 831 1066 842 1071
rect -76 945 -71 950
rect 165 945 170 950
rect 309 915 326 920
rect 837 916 841 921
rect 837 895 842 916
rect 1014 907 1017 912
rect 831 890 842 895
rect -76 769 -71 774
rect 165 769 170 774
rect 309 739 326 744
rect 837 740 841 745
rect 837 719 842 740
rect 831 714 842 719
rect 920 612 925 617
rect -76 593 -71 598
rect 165 593 170 598
rect 309 563 326 568
rect 837 564 841 569
rect 837 543 842 564
rect 831 538 842 543
<< m2contact >>
rect 198 1856 203 1861
rect -71 1825 -66 1830
rect 160 1825 165 1830
rect 198 1795 203 1800
rect 385 1793 390 1798
rect 646 1796 651 1801
rect 900 1793 905 1798
rect 198 1680 203 1685
rect -71 1649 -66 1654
rect 160 1649 165 1654
rect 198 1619 203 1624
rect 385 1617 390 1622
rect 646 1620 651 1625
rect 900 1617 905 1622
rect 198 1504 203 1509
rect -71 1473 -66 1478
rect 160 1473 165 1478
rect 198 1443 203 1448
rect 385 1441 390 1446
rect 646 1444 651 1449
rect 900 1441 905 1446
rect 198 1328 203 1333
rect -71 1297 -66 1302
rect 160 1297 165 1302
rect 198 1267 203 1272
rect 385 1265 390 1270
rect 646 1268 651 1273
rect 900 1265 905 1270
rect 198 1152 203 1157
rect -71 1121 -66 1126
rect 160 1121 165 1126
rect 198 1091 203 1096
rect 385 1089 390 1094
rect 646 1092 651 1097
rect 900 1089 905 1094
rect 198 976 203 981
rect -71 945 -66 950
rect 160 945 165 950
rect 198 915 203 920
rect 385 913 390 918
rect 646 916 651 921
rect 900 913 905 918
rect 1017 907 1022 912
rect 198 800 203 805
rect -71 769 -66 774
rect 160 769 165 774
rect 198 739 203 744
rect 385 737 390 742
rect 646 740 651 745
rect 900 737 905 742
rect 198 624 203 629
rect 915 612 920 617
rect -71 593 -66 598
rect 160 593 165 598
rect 198 563 203 568
rect 385 561 390 566
rect 646 564 651 569
rect 900 561 905 566
<< pm12contact >>
rect 477 1874 482 1879
rect 425 1801 430 1806
rect 587 1801 592 1806
rect 477 1698 482 1703
rect 425 1625 430 1630
rect 587 1625 592 1630
rect 477 1522 482 1527
rect 425 1449 430 1454
rect 587 1449 592 1454
rect 477 1346 482 1351
rect 425 1273 430 1278
rect 587 1273 592 1278
rect 477 1170 482 1175
rect 425 1097 430 1102
rect 587 1097 592 1102
rect 477 994 482 999
rect 425 921 430 926
rect 587 921 592 926
rect 477 818 482 823
rect 425 745 430 750
rect 587 745 592 750
rect 477 642 482 647
rect 425 569 430 574
rect 587 569 592 574
<< metal2 >>
rect 1012 893 1017 898
rect 582 569 587 574
<< m234contact >>
rect 472 1874 477 1879
rect 193 1856 198 1861
rect -76 1825 -71 1830
rect 165 1825 170 1830
rect 430 1801 435 1806
rect 193 1795 198 1800
rect 390 1793 395 1798
rect 651 1796 656 1801
rect 905 1793 910 1798
rect 472 1698 477 1703
rect 193 1680 198 1685
rect -76 1649 -71 1654
rect 165 1649 170 1654
rect 430 1625 435 1630
rect 193 1619 198 1624
rect 390 1617 395 1622
rect 651 1620 656 1625
rect 905 1617 910 1622
rect 472 1522 477 1527
rect 193 1504 198 1509
rect -76 1473 -71 1478
rect 165 1473 170 1478
rect 430 1449 435 1454
rect 193 1443 198 1448
rect 390 1441 395 1446
rect 651 1444 656 1449
rect 905 1441 910 1446
rect 472 1346 477 1351
rect 193 1328 198 1333
rect -76 1297 -71 1302
rect 165 1297 170 1302
rect 430 1273 435 1278
rect 193 1267 198 1272
rect 390 1265 395 1270
rect 651 1268 656 1273
rect 905 1265 910 1270
rect 472 1170 477 1175
rect 193 1152 198 1157
rect -76 1121 -71 1126
rect 165 1121 170 1126
rect 430 1097 435 1102
rect 193 1091 198 1096
rect 390 1089 395 1094
rect 651 1092 656 1097
rect 905 1089 910 1094
rect 472 994 477 999
rect 193 976 198 981
rect -76 945 -71 950
rect 165 945 170 950
rect 430 921 435 926
rect 193 915 198 920
rect 390 913 395 918
rect 651 916 656 921
rect 905 913 910 918
rect 1017 912 1022 917
rect 1017 893 1022 898
rect 472 818 477 823
rect 193 800 198 805
rect -76 769 -71 774
rect 165 769 170 774
rect 430 745 435 750
rect 193 739 198 744
rect 390 737 395 742
rect 651 740 656 745
rect 905 737 910 742
rect 472 642 477 647
rect 193 624 198 629
rect 915 607 920 612
rect -76 593 -71 598
rect 165 593 170 598
rect 430 569 435 574
rect 193 563 198 568
rect 390 561 395 566
rect 651 564 656 569
rect 905 561 910 566
use latch  latch_4
timestamp 1765416915
transform -1 0 -351 0 1 463
box -392 82 -333 1369
use staticizer  staticizer_1
timestamp 1765334200
transform -1 0 43 0 1 1753
box 61 -1215 120 78
use latch  latch_0
timestamp 1765416915
transform 1 0 445 0 1 463
box -392 82 -333 1369
use staticizer  staticizer_0
timestamp 1765334200
transform 1 0 51 0 1 1753
box 61 -1215 120 78
use latch  latch_2
timestamp 1765416915
transform 1 0 982 0 1 459
box -392 82 -333 1369
use shift  shift_0
timestamp 1765416915
transform 1 0 798 0 1 2153
box -138 -1615 46 -268
use addsub  addsub_0
timestamp 1765338694
transform 1 0 421 0 1 712
box -14 -174 166 1225
use latch  latch_1
timestamp 1765416915
transform 1 0 721 0 1 456
box -392 82 -333 1369
use fblock  fblock_0
timestamp 1765416915
transform 1 0 281 0 1 2993
box -80 -2455 50 -1047
use reg  reg_0
timestamp 1765316199
transform 1 0 938 0 1 936
box -14 -398 76 940
use latch  latch_3
timestamp 1765416915
transform 1 0 1236 0 1 456
box -392 82 -333 1369
<< end >>
