magic
tech scmos
timestamp 1765746500
<< metal1 >>
rect -14 908 1 913
rect 75 846 76 851
rect 75 837 76 842
rect -14 732 1 737
rect 75 670 76 675
rect 75 661 76 666
rect -14 556 1 561
rect 75 494 76 499
rect 75 485 76 490
rect -14 380 1 385
rect 75 318 76 323
rect 75 309 76 314
rect -14 204 1 209
rect 75 142 76 147
rect 75 133 76 138
rect -14 28 1 33
rect 75 -34 76 -29
rect 75 -43 76 -38
rect -14 -148 1 -143
rect 75 -210 76 -205
rect 75 -219 76 -214
rect -14 -324 1 -319
rect 75 -386 76 -381
rect 75 -395 76 -390
<< metal2 >>
rect -14 -398 -9 940
<< metal3 >>
rect -3 -398 2 940
rect 6 -398 11 940
rect 24 -398 29 940
rect 70 -398 75 940
use reg_one  reg_one_4
timestamp 1765746319
transform 1 0 2 0 1 331
box -11 -27 74 81
use reg_one  reg_one_6
timestamp 1765746319
transform 1 0 2 0 1 683
box -11 -27 74 81
use reg_one  reg_one_7
timestamp 1765746319
transform 1 0 2 0 1 859
box -11 -27 74 81
use reg_one  reg_one_5
timestamp 1765746319
transform 1 0 2 0 1 507
box -11 -27 74 81
use reg_one  reg_one_3
timestamp 1765746319
transform 1 0 2 0 1 155
box -11 -27 74 81
use reg_one  reg_one_1
timestamp 1765746319
transform 1 0 2 0 1 -197
box -11 -27 74 81
use reg_one  reg_one_2
timestamp 1765746319
transform 1 0 2 0 1 -21
box -11 -27 74 81
use reg_one  reg_one_0
timestamp 1765746319
transform 1 0 2 0 1 -373
box -11 -27 74 81
<< labels >>
rlabel metal1 75 142 76 147 7 port40
rlabel metal1 75 133 76 138 7 port41
rlabel metal1 -2 204 1 209 3 in4
rlabel metal1 75 318 76 323 7 port30
rlabel metal1 75 309 76 314 7 port31
rlabel metal1 -2 380 1 385 3 in3
rlabel metal1 75 494 76 499 7 port20
rlabel metal1 75 485 76 490 7 port21
rlabel metal1 -2 556 1 561 3 in2
rlabel metal1 75 670 76 675 7 port10
rlabel metal1 75 661 76 666 7 port11
rlabel metal1 -2 732 1 737 3 in1
rlabel metal1 75 846 76 851 7 port00
rlabel metal1 75 837 76 842 7 port01
rlabel metal3 6 935 11 940 5 Vdd!
rlabel metal3 24 935 29 940 5 GND!
rlabel metal1 -2 908 1 913 3 in0
rlabel metal3 70 935 75 940 6 w
rlabel metal3 -3 935 2 940 5 r1
rlabel metal2 -14 935 -9 940 4 r0
rlabel metal1 75 -386 76 -381 7 port70
rlabel metal1 75 -395 76 -390 7 port71
rlabel metal1 -2 -324 1 -319 3 in7
rlabel metal1 75 -210 76 -205 7 port60
rlabel metal1 75 -219 76 -214 7 port61
rlabel metal1 -2 -148 1 -143 3 in6
rlabel metal1 75 -34 76 -29 7 port50
rlabel metal1 75 -43 76 -38 7 port51
rlabel metal1 -2 28 1 33 3 in5
<< end >>
