magic
tech scmos
timestamp 1765767571
<< metal5 >>
rect 10 36 14 40
rect 26 36 30 40
rect 10 32 18 36
rect 22 32 30 36
rect 10 28 30 32
rect 10 10 14 28
rect 18 24 22 28
rect 26 10 30 28
rect 34 36 56 40
rect 34 27 38 36
rect 34 23 56 27
rect 34 14 38 23
rect 60 14 64 40
rect 82 36 86 40
rect 82 32 90 36
rect 82 28 94 32
rect 34 10 56 14
rect 60 10 78 14
rect 82 10 86 28
rect 90 26 95 28
rect 90 24 96 26
rect 91 22 96 24
rect 100 22 104 40
rect 108 36 112 40
rect 124 36 128 40
rect 108 32 116 36
rect 120 32 128 36
rect 132 36 150 40
rect 112 28 124 32
rect 92 18 104 22
rect 96 14 104 18
rect 100 10 104 14
rect 116 10 120 28
rect 132 14 136 36
rect 154 28 158 40
rect 168 28 172 40
rect 154 24 172 28
rect 132 10 150 14
rect 154 10 158 24
rect 168 10 172 24
rect 176 14 180 40
rect 194 14 198 40
rect 176 10 198 14
rect 202 27 206 40
rect 218 35 222 40
rect 214 31 222 35
rect 210 27 218 31
rect 202 23 214 27
rect 202 10 206 23
rect 210 19 218 23
rect 214 15 222 19
rect 218 10 222 15
<< end >>
