magic
tech scmos
timestamp 1765669792
<< nwell >>
rect 72 18 134 47
<< pwell >>
rect 101 17 134 18
rect 72 -7 134 17
<< ntransistor >>
rect 84 6 86 11
rect 93 6 95 11
rect 102 6 104 11
rect 111 6 113 11
rect 120 6 122 11
<< ptransistor >>
rect 84 24 86 34
rect 93 24 95 34
rect 102 24 104 34
rect 111 24 113 34
rect 120 24 122 34
<< ndiffusion >>
rect 83 6 84 11
rect 86 6 87 11
rect 92 6 93 11
rect 95 6 96 11
rect 101 6 102 11
rect 104 6 105 11
rect 110 6 111 11
rect 113 6 114 11
rect 119 6 120 11
rect 122 6 123 11
<< pdiffusion >>
rect 83 24 84 34
rect 86 24 93 34
rect 95 24 102 34
rect 104 24 111 34
rect 113 24 120 34
rect 122 24 123 34
<< ndcontact >>
rect 78 6 83 11
rect 87 6 92 11
rect 96 6 101 11
rect 105 6 110 11
rect 114 6 119 11
rect 123 6 128 11
<< pdcontact >>
rect 78 24 83 34
rect 123 24 128 34
<< psubstratepcontact >>
rect 78 -4 83 1
rect 123 -4 128 1
<< nsubstratencontact >>
rect 78 39 83 44
rect 123 39 128 44
<< polysilicon >>
rect 84 34 86 37
rect 93 34 95 37
rect 102 34 104 37
rect 111 34 113 37
rect 120 34 122 37
rect 84 11 86 24
rect 93 11 95 24
rect 102 11 104 24
rect 111 11 113 24
rect 120 11 122 24
rect 84 3 86 6
rect 93 3 95 6
rect 102 3 104 6
rect 111 3 113 6
rect 120 3 122 6
<< metal1 >>
rect 83 39 123 44
rect 128 39 134 44
rect 78 34 83 39
rect 123 20 128 24
rect 87 15 134 20
rect 87 11 92 15
rect 105 11 110 15
rect 123 11 128 15
rect 78 1 83 6
rect 96 1 101 6
rect 114 1 119 6
rect 83 -4 123 1
rect 128 -4 134 1
<< labels >>
rlabel polysilicon 84 35 86 37 1 a
rlabel polysilicon 93 35 95 37 1 b
rlabel polysilicon 102 35 104 37 1 c
rlabel metal1 129 -4 134 1 7 GND!
rlabel polysilicon 111 35 113 37 1 d
rlabel polysilicon 120 35 122 37 1 e
rlabel metal1 129 39 134 44 7 Vdd!
rlabel metal1 129 15 134 20 7 out
<< end >>
