magic
tech scmos
timestamp 1761285742
<< nwell >>
rect 68 15 135 80
<< pwell >>
rect 68 -24 135 15
<< ntransistor >>
rect 85 -11 87 9
rect 95 -11 97 9
rect 105 -11 107 9
rect 116 -11 118 9
<< ptransistor >>
rect 85 24 87 64
rect 95 24 97 64
rect 105 24 107 64
rect 116 24 118 64
<< ndiffusion >>
rect 79 -11 85 9
rect 87 -11 89 9
rect 94 -11 95 9
rect 97 -11 99 9
rect 104 -11 105 9
rect 107 -11 109 9
rect 114 -11 116 9
rect 118 -11 124 9
<< pdiffusion >>
rect 79 24 85 64
rect 87 24 95 64
rect 97 24 105 64
rect 107 24 116 64
rect 118 24 124 64
<< ndcontact >>
rect 74 -11 79 9
rect 89 -11 94 9
rect 99 -11 104 9
rect 109 -11 114 9
rect 124 -11 129 9
<< pdcontact >>
rect 74 24 79 64
rect 124 24 129 64
<< psubstratepcontact >>
rect 99 -21 104 -16
<< nsubstratencontact >>
rect 99 69 104 74
<< polysilicon >>
rect 85 64 87 67
rect 95 64 97 67
rect 105 64 107 67
rect 116 64 118 67
rect 85 9 87 24
rect 95 9 97 24
rect 105 9 107 24
rect 116 9 118 24
rect 85 -14 87 -11
rect 95 -14 97 -11
rect 105 -14 107 -11
rect 116 -14 118 -11
<< metal1 >>
rect 74 69 99 74
rect 104 69 135 74
rect 74 64 79 69
rect 124 19 129 24
rect 89 14 135 19
rect 89 9 94 14
rect 109 9 114 14
rect 74 -16 79 -11
rect 99 -16 104 -11
rect 124 -16 129 -11
rect 74 -21 99 -16
rect 104 -21 135 -16
<< labels >>
rlabel polysilicon 85 65 87 67 1 a
rlabel polysilicon 95 65 97 67 1 b
rlabel polysilicon 105 65 107 67 1 c
rlabel polysilicon 116 65 118 67 1 d
rlabel metal1 130 69 135 74 7 Vdd!
rlabel metal1 130 14 135 19 7 out
rlabel metal1 130 -21 135 -16 7 GND!
<< end >>
