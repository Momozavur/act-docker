magic
tech scmos
timestamp 1765788557
<< pwell >>
rect 1489 1638 1494 1643
rect 1234 1616 1235 1625
<< polysilicon >>
rect 1684 3210 1686 3223
rect 1611 3198 1669 3200
rect 1621 3187 1669 3189
rect 1631 3176 1669 3178
rect 1684 3043 1686 3046
rect 1656 2983 1657 2985
rect 1655 2958 1657 2983
rect 1683 2969 1685 2981
rect 1655 2956 1669 2958
rect 1298 1802 1300 1815
rect 1309 1802 1311 1815
<< polycontact >>
rect 1684 3223 1689 3228
rect 1606 3198 1611 3203
rect 1616 3187 1621 3192
rect 1626 3176 1631 3181
rect 1685 3162 1690 3167
rect 1684 3102 1689 3107
rect 1681 3046 1686 3051
rect 1651 2983 1656 2988
rect 1681 2981 1686 2986
rect 1832 1790 1837 1795
rect 2332 1790 2337 1795
<< metal1 >>
rect 2644 3285 2649 3286
rect 1331 3254 1336 3259
rect 1663 3217 1668 3227
rect 1705 3217 1710 3227
rect 1662 3158 1667 3168
rect 1685 3167 1690 3169
rect 1706 3160 1711 3168
rect 1711 3149 1721 3154
rect 2460 3134 2465 3139
rect 1649 3125 1667 3130
rect 1649 3089 1655 3125
rect 1682 3102 1684 3107
rect 1649 3084 1665 3089
rect 2470 3087 2475 3092
rect 1664 3047 1669 3066
rect 1661 3042 1669 3047
rect 1474 2925 1479 2930
rect 1474 2861 1479 2866
rect 1474 2797 1479 2802
rect 1679 2796 1684 2925
rect 1474 2733 1479 2738
rect 2308 2704 2317 2713
rect 455 2263 464 2704
rect 455 2244 464 2254
rect 569 2262 578 2704
rect 569 2244 578 2253
rect 683 2263 692 2704
rect 683 2245 692 2254
rect 797 2263 806 2704
rect 797 2245 806 2254
rect 911 2263 920 2704
rect 911 2245 920 2254
rect 1025 2263 1034 2704
rect 1025 2245 1034 2254
rect 1139 2263 1148 2704
rect 1139 2245 1148 2254
rect 1253 2263 1262 2704
rect 2380 2595 2385 2600
rect 2360 2546 2365 2551
rect 1253 2245 1262 2254
rect 2608 2257 2617 2266
rect 2608 2248 2660 2257
rect 1253 1758 1258 1784
rect 1805 1769 1814 1774
rect 2305 1769 2316 1774
rect 1253 1753 1278 1758
rect 1273 1634 1278 1753
rect 1286 1727 1291 1762
rect 1805 1729 1810 1769
rect 1805 1724 1816 1729
rect 1835 1725 1840 1732
rect 2305 1729 2310 1769
rect 2609 1737 2618 1764
rect 2305 1724 2316 1729
rect 2335 1722 2340 1737
rect 2609 1732 2640 1737
rect 2651 1732 2660 2248
rect 2611 1729 2616 1732
rect 2653 1728 2658 1732
rect 351 1561 356 1566
rect 3130 1535 3135 1540
rect 3254 1535 3259 1540
rect 351 1385 356 1390
rect 3130 1359 3135 1364
rect 3254 1359 3259 1364
rect 351 1209 356 1214
rect 3130 1183 3135 1188
rect 3254 1183 3259 1188
rect 351 1033 356 1038
rect 3130 1007 3135 1012
rect 3254 1007 3259 1012
rect 351 857 356 862
rect 3130 831 3135 836
rect 3254 831 3259 836
rect 351 681 356 686
rect 3130 655 3135 660
rect 3254 655 3259 660
rect 351 505 356 510
rect 3130 479 3135 484
rect 3254 479 3259 484
rect 351 329 356 334
rect 3130 303 3135 308
rect 3254 303 3259 308
<< m2contact >>
rect 1596 3253 1601 3258
rect 1684 3253 1689 3258
rect 1705 3096 1710 3101
rect 1666 3007 1671 3012
rect 1667 2975 1672 2980
rect 1351 2896 1360 2905
rect 1351 2832 1360 2841
rect 1679 2791 1684 2796
rect 2344 2786 2353 2795
rect 1351 2768 1360 2777
rect 1351 2704 1360 2713
rect 2317 2704 2326 2713
rect 2608 2266 2617 2275
rect 1317 1799 1322 1804
rect 2609 1764 2618 1773
rect 1853 1716 1858 1721
rect 1489 1638 1494 1643
rect 1959 1523 1964 1528
rect 1959 1347 1964 1352
rect 1959 1171 1964 1176
rect 1959 995 1964 1000
rect 1959 819 1964 824
rect 1959 643 1964 648
rect 1959 467 1964 472
rect 1959 291 1964 296
<< pm12contact >>
rect 1296 1815 1301 1820
rect 1309 1815 1314 1820
<< metal2 >>
rect 340 3259 345 3262
rect 448 3259 453 3262
rect 603 3259 608 3262
rect 749 3259 754 3262
rect 1601 3253 1684 3258
rect 1671 3007 1674 3012
rect 1669 2980 1674 3007
rect 1672 2975 1674 2980
rect 1705 2972 1710 3096
rect 528 2800 533 2803
rect 642 2800 647 2803
rect 756 2799 761 2802
rect 870 2800 875 2803
rect 984 2800 989 2803
rect 1212 2799 1217 2802
rect 1326 2799 1331 2802
rect 1098 2785 1103 2788
rect 2598 2225 2603 2232
rect 1317 1754 1322 1799
rect 1848 1770 1862 1775
rect 2348 1770 2362 1775
rect 2594 1773 2603 2225
rect 1848 1716 1853 1770
rect 2348 1716 2353 1770
rect 2594 1764 2609 1773
rect 2681 1764 2690 2214
rect 2699 2205 2708 2222
rect 2699 1764 2708 2196
rect 2717 2187 2726 2222
rect 2717 1764 2726 2178
rect 2735 2169 2744 2222
rect 2735 1764 2744 2160
rect 2763 2151 2772 2222
rect 2763 1764 2772 2142
rect 2781 2133 2790 2222
rect 2781 1764 2790 2124
rect 2799 2115 2808 2222
rect 2799 1764 2808 2106
rect 2817 2097 2826 2222
rect 2817 1764 2826 2088
rect 2845 2079 2854 2222
rect 2845 1764 2854 2070
rect 2863 2061 2872 2222
rect 2863 1764 2872 2052
rect 2881 2043 2890 2222
rect 2881 1764 2890 2034
rect 2899 2025 2908 2222
rect 2899 1764 2908 2016
rect 2927 2007 2936 2222
rect 2927 1764 2936 1998
rect 2945 1989 2954 2222
rect 2945 1764 2954 1980
rect 2963 1971 2972 2222
rect 2963 1764 2972 1962
rect 2981 1953 2990 2222
rect 2981 1764 2990 1944
rect 3009 1935 3018 2222
rect 3009 1755 3018 1926
rect 3027 1917 3036 2222
rect 3027 1765 3036 1908
rect 3045 1899 3054 2222
rect 2384 1746 3018 1755
rect 3045 1737 3054 1890
rect 3063 1881 3072 2222
rect 3063 1764 3072 1872
rect 3091 1863 3100 2222
rect 3091 1764 3100 1854
rect 3109 1845 3118 2222
rect 3109 1764 3118 1836
rect 3127 1827 3136 2222
rect 3127 1764 3136 1818
rect 3145 1809 3154 2222
rect 3145 1764 3154 1800
rect 3173 1791 3182 2222
rect 3173 1764 3182 1782
rect 3189 1773 3198 2222
rect 3209 1764 3218 2222
rect 3227 1764 3236 2222
rect 3000 1728 3054 1737
rect 3000 1697 3009 1728
rect 2364 1688 3009 1697
rect 715 1612 782 1617
rect 1452 1612 1457 1616
rect 1559 1612 1564 1616
rect 1666 1612 1671 1616
rect 2364 1617 2373 1688
rect 1866 1612 1871 1615
rect 2366 1615 2373 1617
rect 2366 1612 2371 1615
rect 2473 1612 2478 1616
rect 2666 1612 2671 1616
rect 804 1611 864 1612
rect 804 1607 859 1611
rect 2661 1607 2671 1612
rect 3000 1608 3009 1688
<< m3contact >>
rect 1582 2967 1587 2972
rect 2681 2214 2690 2223
rect 2699 2196 2708 2205
rect 2717 2178 2726 2187
rect 2735 2160 2744 2169
rect 2763 2142 2772 2151
rect 2781 2124 2790 2133
rect 2799 2106 2808 2115
rect 2817 2088 2826 2097
rect 2845 2070 2854 2079
rect 2863 2052 2872 2061
rect 2881 2034 2890 2043
rect 2899 2016 2908 2025
rect 2927 1998 2936 2007
rect 2945 1980 2954 1989
rect 2963 1962 2972 1971
rect 2981 1944 2990 1953
rect 3009 1926 3018 1935
rect 3027 1908 3036 1917
rect 3045 1890 3054 1899
rect 2375 1746 2384 1755
rect 3063 1872 3072 1881
rect 3091 1854 3100 1863
rect 3109 1836 3118 1845
rect 3127 1818 3136 1827
rect 3145 1800 3154 1809
rect 3173 1782 3182 1791
rect 3189 1764 3198 1773
rect 1559 1616 1564 1621
rect 1666 1616 1671 1621
<< m123contact >>
rect 2591 3285 2597 3291
rect 2644 3286 2649 3291
rect 1714 3128 1719 3133
rect 1738 3128 1743 3133
rect 1717 3107 1722 3112
rect 1663 3089 1668 3094
rect 1651 3075 1656 3080
rect 1646 2983 1651 2988
rect 1705 2967 1710 2972
rect 1663 2948 1668 2953
rect 2367 2883 2376 2892
rect 455 2254 464 2263
rect 569 2253 578 2262
rect 683 2254 692 2263
rect 797 2254 806 2263
rect 911 2254 920 2263
rect 1025 2254 1034 2263
rect 1139 2254 1148 2263
rect 1253 2254 1262 2263
rect 1832 1795 1837 1800
rect 2332 1795 2337 1800
rect 3002 1603 3007 1608
rect 1083 1563 1092 1572
<< metal3 >>
rect 1640 2993 1645 3309
rect 1679 3133 1684 3291
rect 2597 3285 2600 3291
rect 1679 3128 1714 3133
rect 1679 3111 1684 3128
rect 1665 3106 1684 3111
rect 1717 3094 1722 3107
rect 1668 3089 1722 3094
rect 1738 3080 1743 3128
rect 1656 3075 1743 3080
rect 1640 2988 1661 2993
rect 1587 2967 1705 2972
rect 1568 2962 1577 2965
rect 1568 2953 2416 2962
rect 1587 2902 2317 2911
rect 2308 2892 2317 2902
rect 2308 2883 2367 2892
rect 2407 2859 2416 2953
rect 1336 2791 1339 2796
rect 2591 2242 2600 3285
rect 1863 2232 2352 2242
rect 2363 2232 2600 2242
rect 411 2196 2699 2205
rect 411 1601 420 2196
rect 453 2195 483 2196
rect 532 2178 2717 2187
rect 532 1576 541 2178
rect 885 2160 2735 2169
rect 885 1684 894 2160
rect 917 2142 2763 2151
rect 917 1684 926 2142
rect 951 2124 2781 2133
rect 951 1684 960 2124
rect 1057 2106 2799 2115
rect 1057 1706 1066 2106
rect 1083 2088 2817 2097
rect 986 1684 991 1689
rect 986 1653 991 1662
rect 715 1621 720 1626
rect 777 1621 782 1626
rect 936 1574 941 1653
rect 1083 1572 1092 2088
rect 1205 2070 2845 2079
rect 1205 1815 1214 2070
rect 1205 1634 1214 1810
rect 1225 2052 2863 2061
rect 1205 1625 1207 1634
rect 1225 1625 1234 2052
rect 1403 2034 2881 2043
rect 1403 1625 1412 2034
rect 1488 2016 2899 2025
rect 1488 1741 1497 2016
rect 1512 1998 2927 2007
rect 1512 1625 1521 1998
rect 1356 1616 1388 1621
rect 1403 1616 1436 1625
rect 1461 1616 1521 1625
rect 1534 1980 2945 1989
rect 1534 1616 1543 1980
rect 1641 1962 2963 1971
rect 1564 1616 1602 1621
rect 1641 1616 1650 1962
rect 1671 1616 1709 1621
rect 1748 1616 1757 1962
rect 1830 1944 2981 1953
rect 1830 1800 1842 1944
rect 1875 1926 3009 1935
rect 1875 1620 1884 1926
rect 1948 1908 3027 1917
rect 1429 1612 1434 1616
rect 1463 1612 1468 1616
rect 1536 1612 1541 1616
rect 1570 1612 1575 1616
rect 1597 1612 1602 1616
rect 1643 1612 1648 1616
rect 1677 1612 1682 1616
rect 1704 1611 1709 1616
rect 1750 1612 1755 1616
rect 1877 1615 1882 1620
rect 1948 1615 1957 1908
rect 2200 1890 3045 1899
rect 2200 1622 2209 1890
rect 2330 1872 3063 1881
rect 2330 1800 2342 1872
rect 2448 1854 3091 1863
rect 1950 1612 1955 1615
rect 2375 1620 2384 1746
rect 2200 1608 2209 1613
rect 2377 1612 2382 1620
rect 2448 1615 2457 1854
rect 2482 1836 3109 1845
rect 2482 1616 2491 1836
rect 2555 1818 3127 1827
rect 2555 1616 2564 1818
rect 2675 1800 3145 1809
rect 2675 1616 2684 1800
rect 2748 1782 3173 1791
rect 2748 1616 2757 1782
rect 3124 1764 3189 1773
rect 3198 1764 3258 1773
rect 2450 1612 2455 1615
rect 2484 1612 2489 1616
rect 2557 1612 2562 1616
rect 2677 1612 2682 1616
rect 2750 1612 2755 1616
rect 3124 1608 3133 1764
rect 3248 1608 3258 1764
rect 411 1568 416 1571
rect 536 1568 541 1571
rect 859 1561 864 1566
rect 1066 1561 1071 1566
rect 1327 1564 1332 1569
rect 2202 1568 2207 1574
rect 3002 1570 3007 1574
rect 3126 1571 3131 1575
rect 3250 1569 3255 1573
<< m234contact >>
rect 1360 2896 1369 2905
rect 2475 2896 2485 2905
rect 1360 2832 1369 2841
rect 2451 2832 2460 2841
rect 1674 2791 1679 2796
rect 2344 2777 2353 2786
rect 1360 2768 1369 2777
rect 1360 2704 1369 2713
rect 2308 2704 2317 2713
rect 859 1606 864 1611
rect 878 1592 883 1597
rect 1296 1820 1301 1825
rect 1309 1810 1314 1815
rect 1465 1635 1470 1640
rect 1343 1616 1352 1625
rect 1866 1615 1871 1620
rect 1452 1605 1457 1610
rect 1490 1605 1495 1610
rect 2473 1607 2478 1612
rect 478 1546 483 1551
rect 878 1416 883 1421
rect 478 1370 483 1375
rect 878 1240 883 1245
rect 478 1194 483 1199
rect 878 1064 883 1069
rect 478 1018 483 1023
rect 878 888 883 893
rect 478 842 483 847
rect 878 712 883 717
rect 478 666 483 671
rect 878 536 883 541
rect 478 490 483 495
rect 878 360 883 365
rect 478 314 483 319
<< m4contact >>
rect 1640 3309 1645 3314
rect 1679 3291 1684 3296
rect 2591 3291 2600 3300
rect 2642 3291 2651 3300
rect 1413 2955 1422 2964
rect 1531 2955 1540 2964
rect 1339 2791 1344 2796
rect 1852 2232 1863 2242
rect 2352 2232 2363 2242
rect 936 1653 941 1658
rect 981 1653 986 1658
rect 1205 1810 1214 1815
rect 1207 1625 1216 1634
rect 1225 1616 1234 1625
rect 1857 1738 1862 1743
rect 2357 1738 2362 1743
rect 2200 1613 2209 1622
rect 2511 1607 2516 1612
rect 469 1506 474 1511
rect 469 1330 474 1335
rect 469 1154 474 1159
rect 469 978 474 983
rect 469 802 474 807
rect 469 626 474 631
rect 469 450 474 455
rect 469 274 474 279
<< metal4 >>
rect 1413 3314 2651 3318
rect 1413 3309 1640 3314
rect 1645 3309 2651 3314
rect 1413 2964 1422 3309
rect 2642 3300 2651 3309
rect 1531 3296 2591 3300
rect 1531 3291 1679 3296
rect 1684 3291 2591 3296
rect 1531 2964 1540 3291
rect 1369 2896 2475 2905
rect 1369 2832 2451 2841
rect 1344 2791 1674 2796
rect 1369 2768 2353 2777
rect 1369 2704 2308 2713
rect 1301 1820 1470 1825
rect 1214 1810 1309 1815
rect 941 1653 981 1658
rect 1465 1640 1470 1820
rect 1852 1743 1863 2232
rect 2352 1743 2363 2232
rect 1852 1738 1857 1743
rect 1862 1738 1863 1743
rect 1234 1616 1343 1625
rect 1871 1613 2200 1622
rect 1457 1605 1490 1610
rect 2478 1607 2511 1612
<< m345contact >>
rect 455 2244 464 2254
rect 569 2244 578 2253
rect 683 2245 692 2254
rect 797 2245 806 2254
rect 911 2245 920 2254
rect 1025 2245 1034 2254
rect 1139 2245 1148 2254
rect 1253 2245 1262 2254
<< m5contact >>
rect 476 1551 485 1560
rect 476 1375 485 1384
rect 476 1199 485 1208
rect 476 1023 485 1032
rect 476 847 485 856
rect 476 671 485 680
rect 476 495 485 504
rect 476 319 485 328
<< metal5 >>
rect 455 1560 464 2244
rect 455 1551 476 1560
rect 569 1384 578 2244
rect 485 1375 579 1384
rect 683 1208 692 2245
rect 485 1199 692 1208
rect 797 1032 806 2245
rect 485 1023 806 1032
rect 911 856 920 2245
rect 485 847 920 856
rect 1025 680 1034 2245
rect 485 671 1034 680
rect 1139 504 1148 2245
rect 485 495 1148 504
rect 1139 494 1148 495
rect 1253 328 1262 2245
rect 485 319 1262 328
use 2and  2and_0
timestamp 1765747547
transform -1 0 1396 0 1 1729
box 68 29 138 82
use latch_one  latch_one_0
timestamp 1765002978
transform 0 -1 1796 -1 0 1779
box -11 -67 48 -12
use latch_one  latch_one_1
timestamp 1765002978
transform 0 -1 2296 -1 0 1779
box -11 -67 48 -12
use datapath  datapath_0
timestamp 1765779093
transform 1 0 431 0 1 -264
box -81 532 2885 2021
use 2and  2and_1
timestamp 1765747547
transform 0 1 1631 -1 0 3054
box 68 29 138 82
use staticizer_one  staticizer_one_0
timestamp 1765746506
transform 0 1 1717 -1 0 3158
box 54 -61 113 -1
use inv  inv_1
timestamp 1765001281
transform 1 0 1724 0 1 3117
box -10 -13 20 40
use latch_one  latch_one_3
timestamp 1765002978
transform 0 1 1725 -1 0 3034
box -11 -67 48 -12
use inv  inv_0
timestamp 1765001281
transform 0 1 1673 -1 0 3243
box -10 -13 20 40
use 4nor  4nor_0
timestamp 1765673320
transform 0 1 1666 -1 0 3295
box 72 -6 132 47
use latch_one  latch_one_2
timestamp 1765002978
transform 0 1 1726 -1 0 3152
box -11 -67 48 -12
use rom  rom_0
timestamp 1765759847
transform 1 0 2676 0 1 3129
box -350 -907 584 162
use control  control_0
timestamp 1765779093
transform -1 0 1314 0 -1 3151
box -317 -140 974 447
use ring  ring_0
timestamp 1765052771
transform 1 0 179 0 1 3594
box -207 -3603 3499 111
<< labels >>
rlabel metal1 351 1561 356 1566 3 data_out0
rlabel metal1 351 1385 356 1390 3 data_out1
rlabel metal1 351 1209 356 1214 3 data_out2
rlabel metal1 351 1033 356 1038 3 data_out3
rlabel metal1 351 857 356 862 3 data_out4
rlabel metal1 351 681 356 686 3 data_out5
rlabel metal1 351 505 356 510 3 data_out6
rlabel metal1 351 329 356 334 3 data_out7
rlabel m234contact 478 314 483 319 1 data_in7
rlabel m234contact 478 490 483 495 1 data_in6
rlabel m234contact 478 666 483 671 1 data_in5
rlabel m234contact 478 842 483 847 1 data_in4
rlabel m234contact 478 1018 483 1023 1 data_in3
rlabel m234contact 478 1194 483 1199 1 data_in2
rlabel m234contact 478 1370 483 1375 1 data_in1
rlabel metal2 3209 2045 3218 2054 1 r_-w
rlabel metal1 3254 1359 3259 1364 1 addr_out9
rlabel metal1 3254 1535 3259 1540 1 addr_out8
rlabel metal1 3254 1183 3259 1188 1 addr_out10
rlabel metal1 3254 1007 3259 1012 1 addr_out11
rlabel metal1 3254 831 3259 836 1 addr_out12
rlabel metal1 3254 655 3259 660 1 addr_out13
rlabel metal1 3254 479 3259 484 1 addr_out14
rlabel metal1 3254 303 3259 308 1 addr_out15
rlabel metal1 3130 1536 3135 1540 1 addr_out0
rlabel metal1 3130 1360 3135 1364 1 addr_out1
rlabel metal1 3130 1184 3135 1188 1 addr_out2
rlabel metal1 3130 1008 3135 1012 1 addr_out3
rlabel metal1 3130 832 3135 836 1 addr_out4
rlabel metal1 3130 656 3135 660 1 addr_out5
rlabel metal1 3130 480 3135 484 1 addr_out6
rlabel metal1 3130 304 3135 308 1 addr_out7
rlabel metal1 2360 2546 2365 2551 1 s3
rlabel metal1 2380 2595 2385 2600 1 s2
rlabel metal1 2460 3134 2465 3139 1 s1
rlabel metal1 2644 3285 2649 3291 1 phi1
rlabel metal1 2470 3087 2475 3092 1 s0
rlabel metal3 411 1568 416 1571 1 rd_dataout
rlabel metal3 536 1568 541 1571 1 ld_datain
rlabel metal3 715 1621 720 1626 1 os_u
rlabel metal3 777 1621 782 1626 1 os_s
rlabel metal3 859 1561 864 1566 1 ros
rlabel metal3 887 1684 892 1689 1 fb_g3
rlabel metal3 919 1684 924 1689 1 fb_g2
rlabel metal3 953 1684 958 1689 1 fb_g1
rlabel metal3 986 1684 991 1689 1 fb_g0
rlabel metal3 1066 1561 1071 1566 1 rfb
rlabel m123contact 1087 1565 1092 1570 1 as_sub
rlabel metal1 1273 1634 1278 1639 1 as_cin
rlabel m234contact 1345 1616 1350 1621 1 A_r0
rlabel metal3 1356 1616 1361 1621 1 A_r1
rlabel metal3 1327 1564 1332 1569 1 ras
rlabel m234contact 878 1592 883 1597 1 ry0
rlabel m234contact 878 1416 883 1421 1 ry1
rlabel m234contact 878 1240 883 1245 1 ry2
rlabel m234contact 878 1064 883 1069 1 ry3
rlabel m234contact 878 888 883 893 1 ry4
rlabel m234contact 878 712 883 717 1 ry5
rlabel m234contact 878 536 883 541 1 ry6
rlabel m234contact 878 360 883 365 1 ry7
rlabel m4contact 469 1506 474 1511 1 rx0
rlabel m4contact 469 1330 474 1335 1 rx1
rlabel m4contact 469 1154 474 1159 1 rx2
rlabel m4contact 469 978 474 983 1 rx3
rlabel m4contact 469 802 474 807 1 rx4
rlabel m4contact 469 626 474 631 1 rx5
rlabel m4contact 469 450 474 455 1 rx6
rlabel m4contact 469 274 474 279 1 rx7
rlabel m2contact 1959 1523 1964 1526 1 rx_PCL0
rlabel m2contact 1959 1347 1964 1350 1 rx_PCL1
rlabel m2contact 1959 1171 1964 1174 1 rx_PCL2
rlabel m2contact 1959 995 1964 998 1 rx_PCL3
rlabel m2contact 1959 819 1964 822 1 rx_PCL4
rlabel m2contact 1959 643 1964 646 1 rx_PCL5
rlabel m2contact 1959 467 1964 470 1 rx_PCL6
rlabel m2contact 1959 291 1964 294 1 rx_PCL7
rlabel metal3 1429 1612 1434 1616 1 A_w
rlabel metal2 1452 1612 1457 1616 1 DB_r0
rlabel metal3 1463 1612 1468 1616 1 DB_r1
rlabel metal3 1536 1612 1541 1616 1 DB_w
rlabel metal2 1559 1612 1564 1616 1 X_r0
rlabel metal3 1570 1612 1575 1616 1 X_r1
rlabel metal3 1643 1612 1648 1616 1 X_w
rlabel metal2 1666 1612 1671 1616 1 Y_r0
rlabel metal3 1677 1612 1682 1616 1 Y_r1
rlabel metal3 1750 1612 1755 1616 1 Y_w
rlabel metal3 1876 1622 1881 1627 1 PCL_r1
rlabel metal2 1866 1612 1871 1615 1 PCL_r0
rlabel metal3 1950 1612 1955 1615 1 PCL_w
rlabel metal3 2202 1571 2207 1574 1 rPCplus1L
rlabel metal2 2366 1612 2371 1615 1 PCH_r0
rlabel metal3 2377 1612 2382 1615 1 PCH_r1
rlabel metal3 2450 1612 2455 1615 1 PCH_w
rlabel metal2 2473 1612 2478 1616 1 ABL_r0
rlabel metal3 2484 1612 2489 1616 1 ABL_r1
rlabel metal3 2557 1612 2562 1616 1 ABL_w
rlabel metal1 2635 1732 2640 1736 1 ABH_w_sel
rlabel metal2 2666 1612 2671 1616 1 ABH_r0
rlabel metal3 2677 1612 2682 1616 1 ABH_r1
rlabel metal3 2750 1612 2755 1616 1 ABH_w
rlabel metal3 3002 1570 3007 1574 1 rPCplus1H
rlabel metal3 3126 1572 3131 1575 1 rd_addrL
rlabel metal3 3250 1570 3255 1573 1 rd_addrH
rlabel metal1 2335 1729 2339 1732 1 PCH_w_sel
rlabel metal1 1835 1725 1840 1732 1 PCL_w_sel
rlabel m123contact 2591 3285 2596 3291 1 phi0
rlabel metal3 1491 1741 1496 1746 1 Cflag_w
rlabel m2contact 1489 1638 1494 1643 1 Cflag
rlabel space 177 3682 319 3696 1 Vdd!
rlabel space 632 3688 640 3700 1 phi0
rlabel space 982 3690 990 3702 1 phi1
rlabel space 1332 3688 1340 3705 1 reset
rlabel space -29 3452 -17 3460 1 r-w_
rlabel space -29 3102 -17 3110 1 d0
rlabel space -29 2752 -17 2760 1 d1
rlabel space -29 2402 -17 2410 1 d2
rlabel space -29 2052 -17 2060 1 d3
rlabel space -29 1702 -17 1710 1 d4
rlabel space -29 1352 -18 1360 1 d5
rlabel space -29 1002 -17 1010 1 d6
rlabel space -29 652 -17 660 1 d7
rlabel space -28 198 -14 340 1 GND!
rlabel space 558 -9 566 3 1 a15
rlabel space 908 -9 916 3 1 a14
rlabel space 1258 -9 1266 3 1 a13
rlabel space 1608 -9 1616 3 1 a12
rlabel space 1958 -9 1966 3 1 a11
rlabel space 2308 -9 2316 3 1 a10
rlabel space 2658 -9 2666 3 1 a9
rlabel space 3008 -9 3016 3 1 a8
rlabel space 3328 -8 3470 6 1 Vdd!
rlabel space 3665 228 3677 236 1 a7
rlabel space 3665 578 3677 586 1 a6
rlabel space 3665 928 3677 936 1 a5
rlabel space 3665 1278 3677 1286 1 a4
rlabel space 3665 1628 3677 1636 1 a3
rlabel space 3665 1978 3677 1986 1 a2
rlabel space 3665 2328 3677 2336 1 a1
rlabel space 3665 2678 3677 2686 1 a0
rlabel space 3662 3348 3676 3490 1 GND!
rlabel m234contact 478 1546 483 1551 1 data_in0
rlabel metal1 1331 3254 1336 3259 1 rst
rlabel metal2 528 2800 533 2803 1 IR0
rlabel metal2 642 2800 647 2803 1 IR1
rlabel metal2 756 2799 761 2802 1 IR2
rlabel metal2 870 2800 875 2803 1 IR3
rlabel metal2 984 2800 989 2803 1 IR4
rlabel metal2 1098 2785 1103 2788 1 IR5
rlabel metal2 1212 2799 1217 2802 1 IR6
rlabel metal2 1326 2799 1331 2802 1 IR7
rlabel metal2 749 3259 754 3262 1 s0'
rlabel metal2 603 3259 608 3262 1 s1'
rlabel metal2 448 3259 453 3262 1 s2'
rlabel metal1 1474 2925 1479 2930 1 s0_int
rlabel metal1 1474 2861 1479 2866 1 s1_int
rlabel metal1 1474 2797 1479 2802 1 s2_int
rlabel metal1 1474 2733 1479 2738 1 s3_int
rlabel metal2 340 3259 345 3262 1 s3'
rlabel polycontact 1685 3162 1690 3167 1 IR_w_next
rlabel m4contact 1339 2791 1344 2796 1 IR_w
rlabel polycontact 1684 3102 1689 3107 1 IR_w_int
rlabel polycontact 1681 2981 1686 2986 1 IR_w_latched
<< end >>
