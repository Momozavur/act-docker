magic
tech scmos
timestamp 1765311847
<< metal1 >>
rect -80 -1137 -79 -1132
rect -80 -1198 -79 -1193
rect 18 -1198 28 -1193
rect -80 -1313 -79 -1308
rect -80 -1374 -79 -1369
rect 18 -1374 28 -1369
rect -80 -1489 -79 -1484
rect -80 -1550 -79 -1545
rect 18 -1550 28 -1545
rect -80 -1665 -79 -1660
rect -80 -1726 -79 -1721
rect 18 -1726 28 -1721
rect -80 -1841 -79 -1836
rect -80 -1902 -79 -1897
rect 18 -1902 28 -1897
rect -80 -2017 -79 -2012
rect -80 -2078 -79 -2073
rect 18 -2078 28 -2073
rect -80 -2193 -79 -2188
rect -80 -2254 -79 -2249
rect 18 -2254 28 -2249
rect -80 -2369 -79 -2364
rect -80 -2430 -79 -2425
rect 18 -2430 28 -2425
<< m3contact >>
rect -30 -1159 -25 -1154
rect -30 -1335 -25 -1330
rect -30 -1511 -25 -1506
rect -30 -1687 -25 -1682
rect -30 -1863 -25 -1858
rect -30 -2039 -25 -2034
rect -30 -2215 -25 -2210
rect -30 -2391 -25 -2386
<< m123contact >>
rect 42 -1056 47 -1051
rect -79 -1076 -74 -1071
rect -47 -1076 -42 -1071
rect -13 -1076 -8 -1071
rect 20 -1076 25 -1071
rect 42 -1232 47 -1227
rect -79 -1252 -74 -1247
rect -47 -1252 -42 -1247
rect -13 -1252 -8 -1247
rect 20 -1252 25 -1247
rect 42 -1408 47 -1403
rect -79 -1428 -74 -1423
rect -47 -1428 -42 -1423
rect -13 -1428 -8 -1423
rect 20 -1428 25 -1423
rect 42 -1584 47 -1579
rect -79 -1604 -74 -1599
rect -47 -1604 -42 -1599
rect -13 -1604 -8 -1599
rect 20 -1604 25 -1599
rect 42 -1760 47 -1755
rect -79 -1780 -74 -1775
rect -47 -1780 -42 -1775
rect -13 -1780 -8 -1775
rect 20 -1780 25 -1775
rect 42 -1936 47 -1931
rect -79 -1956 -74 -1951
rect -47 -1956 -42 -1951
rect -13 -1956 -8 -1951
rect 20 -1956 25 -1951
rect 42 -2112 47 -2107
rect -79 -2132 -74 -2127
rect -47 -2132 -42 -2127
rect -13 -2132 -8 -2127
rect 20 -2132 25 -2127
rect 42 -2288 47 -2283
rect -79 -2308 -74 -2303
rect -47 -2308 -42 -2303
rect -13 -2308 -8 -2303
rect 20 -2308 25 -2303
<< metal3 >>
rect -79 -1247 -74 -1076
rect -79 -1423 -74 -1252
rect -79 -1599 -74 -1428
rect -79 -1775 -74 -1604
rect -79 -1951 -74 -1780
rect -79 -2127 -74 -1956
rect -79 -2303 -74 -2132
rect -47 -1247 -42 -1076
rect -47 -1423 -42 -1252
rect -47 -1599 -42 -1428
rect -47 -1775 -42 -1604
rect -47 -1951 -42 -1780
rect -47 -2127 -42 -1956
rect -47 -2303 -42 -2132
rect -30 -1330 -25 -1159
rect -30 -1506 -25 -1335
rect -30 -1682 -25 -1511
rect -30 -1858 -25 -1687
rect -30 -2034 -25 -1863
rect -30 -2210 -25 -2039
rect -30 -2386 -25 -2215
rect -13 -1247 -8 -1076
rect -13 -1423 -8 -1252
rect -13 -1599 -8 -1428
rect -13 -1775 -8 -1604
rect -13 -1951 -8 -1780
rect -13 -2127 -8 -1956
rect -13 -2303 -8 -2132
rect 20 -1247 25 -1076
rect 20 -1423 25 -1252
rect 20 -1599 25 -1428
rect 20 -1775 25 -1604
rect 20 -1951 25 -1780
rect 20 -2127 25 -1956
rect 20 -2303 25 -2132
rect 42 -1227 47 -1056
rect 42 -1403 47 -1232
rect 42 -1579 47 -1408
rect 42 -1755 47 -1584
rect 42 -1931 47 -1760
rect 42 -2107 47 -1936
rect 42 -2283 47 -2112
use fblock_one  fblock_one_0
timestamp 1765250278
transform 1 0 -75 0 1 -1133
box -5 -90 125 86
use fblock_one  fblock_one_1
timestamp 1765250278
transform 1 0 -75 0 1 -1309
box -5 -90 125 86
use fblock_one  fblock_one_2
timestamp 1765250278
transform 1 0 -75 0 1 -1485
box -5 -90 125 86
use fblock_one  fblock_one_3
timestamp 1765250278
transform 1 0 -75 0 1 -1661
box -5 -90 125 86
use fblock_one  fblock_one_4
timestamp 1765250278
transform 1 0 -75 0 1 -1837
box -5 -90 125 86
use fblock_one  fblock_one_5
timestamp 1765250278
transform 1 0 -75 0 1 -2013
box -5 -90 125 86
use fblock_one  fblock_one_6
timestamp 1765250278
transform 1 0 -75 0 1 -2189
box -5 -90 125 86
use fblock_one  fblock_one_7
timestamp 1765250278
transform 1 0 -75 0 1 -2365
box -5 -90 125 86
<< labels >>
rlabel m123contact -79 -1076 -74 -1071 3 g3
rlabel m123contact -47 -1076 -42 -1071 1 g2
rlabel m123contact -13 -1076 -8 -1071 1 g1
rlabel m123contact 20 -1076 25 -1071 1 g0
rlabel m123contact 42 -1056 47 -1051 1 Vdd!
rlabel m3contact -30 -1159 -25 -1154 1 GND!
rlabel metal1 -80 -1137 -79 -1132 3 b0
rlabel metal1 -80 -1198 -79 -1193 3 a0
rlabel metal1 -80 -1374 -79 -1369 3 a1
rlabel metal1 -80 -1550 -79 -1545 3 a2
rlabel metal1 -80 -1726 -79 -1721 3 a3
rlabel metal1 -80 -2078 -79 -2073 3 a5
rlabel metal1 -80 -2254 -79 -2249 3 a6
rlabel metal1 -80 -2430 -79 -2425 3 a7
rlabel metal1 -80 -1902 -79 -1897 3 a4
rlabel metal1 -80 -1313 -79 -1308 3 b1
rlabel metal1 -80 -1489 -79 -1484 3 b2
rlabel metal1 -80 -1665 -79 -1660 3 b3
rlabel metal1 -80 -1841 -79 -1836 3 b4
rlabel metal1 -80 -2017 -79 -2012 3 b5
rlabel metal1 -80 -2193 -79 -2188 3 b6
rlabel metal1 -80 -2369 -79 -2364 3 b7
rlabel metal1 25 -1198 28 -1193 1 f0
rlabel metal1 25 -1374 28 -1369 1 f1
rlabel metal1 25 -1550 28 -1545 1 f2
rlabel metal1 25 -1726 28 -1721 1 f3
rlabel metal1 25 -1902 28 -1897 1 f4
rlabel metal1 25 -2078 28 -2073 1 f5
rlabel metal1 25 -2254 28 -2249 1 f6
rlabel metal1 25 -2430 28 -2425 1 f7
<< end >>
