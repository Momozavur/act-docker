magic
tech scmos
timestamp 1765495026
<< polysilicon >>
rect 678 1804 679 1806
rect 678 1628 679 1630
rect 678 1452 679 1454
rect 678 1276 679 1278
rect 678 1100 679 1102
rect 678 924 679 926
rect 678 748 679 750
rect 678 572 679 574
<< polycontact >>
rect -20 1800 -15 1805
rect 109 1800 114 1805
rect 373 1796 378 1801
rect 580 1795 585 1800
rect -20 1624 -15 1629
rect 109 1624 114 1629
rect 373 1620 378 1625
rect 580 1619 585 1624
rect -20 1448 -15 1453
rect 109 1448 114 1453
rect 373 1444 378 1449
rect 580 1443 585 1448
rect -20 1272 -15 1277
rect 109 1272 114 1277
rect 373 1268 378 1273
rect 580 1267 585 1272
rect -20 1096 -15 1101
rect 109 1096 114 1101
rect 373 1092 378 1097
rect 580 1091 585 1096
rect -20 920 -15 925
rect 109 920 114 925
rect 373 916 378 921
rect 580 915 585 920
rect -20 744 -15 749
rect 109 744 114 749
rect 373 740 378 745
rect 580 739 585 744
rect -20 568 -15 573
rect 109 568 114 573
rect 373 564 378 569
rect 580 563 585 568
<< metal1 >>
rect 910 1844 915 1849
rect 1017 1844 1022 1849
rect 1124 1844 1129 1849
rect 1231 1844 1236 1849
rect -76 1825 -71 1830
rect 369 1796 373 1801
rect 369 1775 374 1796
rect 563 1795 580 1800
rect 1004 1787 1007 1792
rect 1111 1787 1114 1792
rect 1218 1787 1221 1792
rect 1325 1787 1328 1792
rect 363 1770 374 1775
rect 910 1668 915 1673
rect 1017 1668 1022 1673
rect 1124 1668 1129 1673
rect 1231 1668 1236 1673
rect -76 1649 -71 1654
rect 369 1620 373 1625
rect 369 1599 374 1620
rect 563 1619 580 1624
rect 1004 1611 1007 1616
rect 1111 1611 1114 1616
rect 1218 1611 1221 1616
rect 1325 1611 1328 1616
rect 363 1594 374 1599
rect 910 1492 915 1497
rect 1017 1492 1022 1497
rect 1124 1492 1129 1497
rect 1231 1492 1236 1497
rect -76 1473 -71 1478
rect 369 1444 373 1449
rect 369 1423 374 1444
rect 563 1443 580 1448
rect 1004 1435 1007 1440
rect 1111 1435 1114 1440
rect 1218 1435 1221 1440
rect 1325 1435 1328 1440
rect 363 1418 374 1423
rect 910 1316 915 1321
rect 1017 1316 1022 1321
rect 1124 1316 1129 1321
rect 1231 1316 1236 1321
rect -76 1297 -71 1302
rect 369 1268 373 1273
rect 369 1247 374 1268
rect 563 1267 580 1272
rect 1004 1259 1007 1264
rect 1111 1259 1114 1264
rect 1218 1259 1221 1264
rect 1325 1259 1328 1264
rect 363 1242 374 1247
rect 910 1140 915 1145
rect 1017 1140 1022 1145
rect 1124 1140 1129 1145
rect 1231 1140 1236 1145
rect -76 1121 -71 1126
rect 369 1092 373 1097
rect 369 1071 374 1092
rect 563 1091 580 1096
rect 1004 1083 1007 1088
rect 1111 1083 1114 1088
rect 1218 1083 1221 1088
rect 1325 1083 1328 1088
rect 363 1066 374 1071
rect 910 964 915 969
rect 1017 964 1022 969
rect 1124 964 1129 969
rect 1231 964 1236 969
rect -76 945 -71 950
rect 369 916 373 921
rect 369 895 374 916
rect 563 915 580 920
rect 1004 907 1007 912
rect 1111 907 1114 912
rect 1218 907 1221 912
rect 1325 907 1328 912
rect 363 890 374 895
rect 910 788 915 793
rect 1017 788 1022 793
rect 1124 788 1129 793
rect 1231 788 1236 793
rect -76 769 -71 774
rect 369 740 373 745
rect 369 719 374 740
rect 563 739 580 744
rect 1004 731 1007 736
rect 1111 731 1114 736
rect 1218 731 1221 736
rect 1325 731 1328 736
rect 363 714 374 719
rect 910 612 915 617
rect 1017 612 1022 617
rect 1124 612 1129 617
rect 1231 612 1236 617
rect -76 593 -71 598
rect 369 564 373 569
rect 369 543 374 564
rect 563 563 580 568
rect 1004 555 1007 560
rect 1111 555 1114 560
rect 1218 555 1221 560
rect 1325 555 1328 560
rect 363 538 374 543
<< m2contact >>
rect 452 1856 457 1861
rect 905 1844 910 1849
rect 1012 1844 1017 1849
rect 1119 1844 1124 1849
rect 1226 1844 1231 1849
rect -71 1825 -66 1830
rect 432 1793 437 1798
rect 452 1795 457 1800
rect 639 1793 644 1798
rect 900 1796 905 1801
rect 1007 1787 1012 1792
rect 1114 1787 1119 1792
rect 1221 1787 1226 1792
rect 1328 1787 1333 1792
rect 452 1680 457 1685
rect 905 1668 910 1673
rect 1012 1668 1017 1673
rect 1119 1668 1124 1673
rect 1226 1668 1231 1673
rect -71 1649 -66 1654
rect 432 1617 437 1622
rect 452 1619 457 1624
rect 639 1617 644 1622
rect 900 1620 905 1625
rect 1007 1611 1012 1616
rect 1114 1611 1119 1616
rect 1221 1611 1226 1616
rect 1328 1611 1333 1616
rect 452 1504 457 1509
rect 905 1492 910 1497
rect 1012 1492 1017 1497
rect 1119 1492 1124 1497
rect 1226 1492 1231 1497
rect -71 1473 -66 1478
rect 432 1441 437 1446
rect 452 1443 457 1448
rect 639 1441 644 1446
rect 900 1444 905 1449
rect 1007 1435 1012 1440
rect 1114 1435 1119 1440
rect 1221 1435 1226 1440
rect 1328 1435 1333 1440
rect 452 1328 457 1333
rect 905 1316 910 1321
rect 1012 1316 1017 1321
rect 1119 1316 1124 1321
rect 1226 1316 1231 1321
rect -71 1297 -66 1302
rect 432 1265 437 1270
rect 452 1267 457 1272
rect 639 1265 644 1270
rect 900 1268 905 1273
rect 1007 1259 1012 1264
rect 1114 1259 1119 1264
rect 1221 1259 1226 1264
rect 1328 1259 1333 1264
rect 452 1152 457 1157
rect 905 1140 910 1145
rect 1012 1140 1017 1145
rect 1119 1140 1124 1145
rect 1226 1140 1231 1145
rect -71 1121 -66 1126
rect 432 1089 437 1094
rect 452 1091 457 1096
rect 639 1089 644 1094
rect 900 1092 905 1097
rect 1007 1083 1012 1088
rect 1114 1083 1119 1088
rect 1221 1083 1226 1088
rect 1328 1083 1333 1088
rect 452 976 457 981
rect 905 964 910 969
rect 1012 964 1017 969
rect 1119 964 1124 969
rect 1226 964 1231 969
rect -71 945 -66 950
rect 432 913 437 918
rect 452 915 457 920
rect 639 913 644 918
rect 900 916 905 921
rect 1007 907 1012 912
rect 1114 907 1119 912
rect 1221 907 1226 912
rect 1328 907 1333 912
rect 452 800 457 805
rect 905 788 910 793
rect 1012 788 1017 793
rect 1119 788 1124 793
rect 1226 788 1231 793
rect -71 769 -66 774
rect 432 737 437 742
rect 452 739 457 744
rect 639 737 644 742
rect 900 740 905 745
rect 1007 731 1012 736
rect 1114 731 1119 736
rect 1221 731 1226 736
rect 1328 731 1333 736
rect 452 624 457 629
rect 905 612 910 617
rect 1012 612 1017 617
rect 1119 612 1124 617
rect 1226 612 1231 617
rect -71 593 -66 598
rect 432 561 437 566
rect 452 563 457 568
rect 639 561 644 566
rect 900 564 905 569
rect 1007 555 1012 560
rect 1114 555 1119 560
rect 1221 555 1226 560
rect 1328 555 1333 560
<< pm12contact >>
rect 731 1874 736 1879
rect 679 1801 684 1806
rect 841 1801 846 1806
rect 731 1698 736 1703
rect 679 1625 684 1630
rect 841 1625 846 1630
rect 731 1522 736 1527
rect 679 1449 684 1454
rect 841 1449 846 1454
rect 731 1346 736 1351
rect 679 1273 684 1278
rect 841 1273 846 1278
rect 731 1170 736 1175
rect 679 1097 684 1102
rect 841 1097 846 1102
rect 731 994 736 999
rect 679 921 684 926
rect 841 921 846 926
rect 731 818 736 823
rect 679 745 684 750
rect 841 745 846 750
rect 731 642 736 647
rect 679 569 684 574
rect 841 569 846 574
<< metal2 >>
rect 447 1795 452 1800
rect 1002 1773 1007 1778
rect 1109 1773 1114 1778
rect 1216 1773 1221 1778
rect 1323 1773 1328 1778
rect 447 1619 452 1624
rect 1002 1597 1007 1602
rect 1109 1597 1114 1602
rect 1216 1597 1221 1602
rect 1323 1597 1328 1602
rect 447 1443 452 1448
rect 1002 1421 1007 1426
rect 1109 1421 1114 1426
rect 1216 1421 1221 1426
rect 1323 1421 1328 1426
rect 447 1267 452 1272
rect 1002 1245 1007 1250
rect 1109 1245 1114 1250
rect 1216 1245 1221 1250
rect 1323 1245 1328 1250
rect 447 1091 452 1096
rect 1002 1069 1007 1074
rect 1109 1069 1114 1074
rect 1216 1069 1221 1074
rect 1323 1069 1328 1074
rect 447 915 452 920
rect 1002 893 1007 898
rect 1109 893 1114 898
rect 1216 893 1221 898
rect 1323 893 1328 898
rect 447 739 452 744
rect 1002 717 1007 722
rect 1109 717 1114 722
rect 1216 717 1221 722
rect 1323 717 1328 722
rect 836 569 841 574
rect 447 563 452 568
rect 1002 541 1007 546
rect 1109 541 1114 546
rect 1216 541 1221 546
rect 1323 541 1328 546
<< m3contact >>
rect 726 1874 731 1879
rect 684 1801 689 1806
rect 726 1698 731 1703
rect 684 1625 689 1630
rect 726 1522 731 1527
rect 684 1449 689 1454
rect 726 1346 731 1351
rect 684 1273 689 1278
rect 726 1170 731 1175
rect 684 1097 689 1102
rect 726 994 731 999
rect 684 921 689 926
rect 726 818 731 823
rect 684 745 689 750
rect 726 642 731 647
rect 684 569 689 574
<< m123contact >>
rect 160 1825 165 1830
rect 160 1649 165 1654
rect 160 1473 165 1478
rect 160 1297 165 1302
rect 160 1121 165 1126
rect 160 945 165 950
rect 160 769 165 774
rect 160 593 165 598
<< metal3 >>
rect 165 1798 170 1830
rect 684 1806 689 1856
rect 447 1775 452 1800
rect 726 1820 731 1874
rect 684 1778 689 1801
rect 905 1801 910 1839
rect 1007 1797 1012 1815
rect 165 1622 170 1654
rect 684 1630 689 1680
rect 447 1599 452 1624
rect 726 1644 731 1698
rect 684 1602 689 1625
rect 905 1625 910 1663
rect 1007 1621 1012 1639
rect 165 1446 170 1478
rect 684 1454 689 1504
rect 447 1423 452 1448
rect 726 1468 731 1522
rect 684 1426 689 1449
rect 905 1449 910 1487
rect 1007 1445 1012 1463
rect 165 1270 170 1302
rect 684 1278 689 1328
rect 447 1247 452 1272
rect 726 1292 731 1346
rect 684 1250 689 1273
rect 905 1273 910 1311
rect 1007 1269 1012 1287
rect 165 1094 170 1126
rect 684 1102 689 1152
rect 447 1071 452 1096
rect 726 1116 731 1170
rect 684 1074 689 1097
rect 905 1097 910 1135
rect 1007 1093 1012 1111
rect 165 918 170 950
rect 684 926 689 976
rect 447 895 452 920
rect 726 940 731 994
rect 684 898 689 921
rect 905 921 910 959
rect 1007 917 1012 935
rect 165 742 170 774
rect 684 750 689 800
rect 447 719 452 744
rect 726 764 731 818
rect 684 722 689 745
rect 905 745 910 783
rect 1007 741 1012 759
rect 165 566 170 598
rect 684 574 689 624
rect 447 543 452 568
rect 726 588 731 642
rect 684 546 689 569
rect 905 569 910 607
rect 1007 565 1012 583
<< m234contact >>
rect 447 1856 452 1861
rect -76 1825 -71 1830
rect 447 1800 452 1805
rect 437 1793 442 1798
rect 905 1839 910 1844
rect 1012 1839 1017 1844
rect 1119 1839 1124 1844
rect 1226 1839 1231 1844
rect 644 1793 649 1798
rect 905 1796 910 1801
rect 1007 1792 1012 1797
rect 1114 1792 1119 1797
rect 1221 1792 1226 1797
rect 1328 1792 1333 1797
rect 1007 1773 1012 1778
rect 1114 1773 1119 1778
rect 1221 1773 1226 1778
rect 1328 1773 1333 1778
rect 447 1680 452 1685
rect -76 1649 -71 1654
rect 447 1624 452 1629
rect 437 1617 442 1622
rect 905 1663 910 1668
rect 1012 1663 1017 1668
rect 1119 1663 1124 1668
rect 1226 1663 1231 1668
rect 644 1617 649 1622
rect 905 1620 910 1625
rect 1007 1616 1012 1621
rect 1114 1616 1119 1621
rect 1221 1616 1226 1621
rect 1328 1616 1333 1621
rect 1007 1597 1012 1602
rect 1114 1597 1119 1602
rect 1221 1597 1226 1602
rect 1328 1597 1333 1602
rect 447 1504 452 1509
rect -76 1473 -71 1478
rect 447 1448 452 1453
rect 437 1441 442 1446
rect 905 1487 910 1492
rect 1012 1487 1017 1492
rect 1119 1487 1124 1492
rect 1226 1487 1231 1492
rect 644 1441 649 1446
rect 905 1444 910 1449
rect 1007 1440 1012 1445
rect 1114 1440 1119 1445
rect 1221 1440 1226 1445
rect 1328 1440 1333 1445
rect 1007 1421 1012 1426
rect 1114 1421 1119 1426
rect 1221 1421 1226 1426
rect 1328 1421 1333 1426
rect 447 1328 452 1333
rect -76 1297 -71 1302
rect 447 1272 452 1277
rect 437 1265 442 1270
rect 905 1311 910 1316
rect 1012 1311 1017 1316
rect 1119 1311 1124 1316
rect 1226 1311 1231 1316
rect 644 1265 649 1270
rect 905 1268 910 1273
rect 1007 1264 1012 1269
rect 1114 1264 1119 1269
rect 1221 1264 1226 1269
rect 1328 1264 1333 1269
rect 1007 1245 1012 1250
rect 1114 1245 1119 1250
rect 1221 1245 1226 1250
rect 1328 1245 1333 1250
rect 447 1152 452 1157
rect -76 1121 -71 1126
rect 447 1096 452 1101
rect 437 1089 442 1094
rect 905 1135 910 1140
rect 1012 1135 1017 1140
rect 1119 1135 1124 1140
rect 1226 1135 1231 1140
rect 644 1089 649 1094
rect 905 1092 910 1097
rect 1007 1088 1012 1093
rect 1114 1088 1119 1093
rect 1221 1088 1226 1093
rect 1328 1088 1333 1093
rect 1007 1069 1012 1074
rect 1114 1069 1119 1074
rect 1221 1069 1226 1074
rect 1328 1069 1333 1074
rect 447 976 452 981
rect -76 945 -71 950
rect 447 920 452 925
rect 437 913 442 918
rect 905 959 910 964
rect 1012 959 1017 964
rect 1119 959 1124 964
rect 1226 959 1231 964
rect 644 913 649 918
rect 905 916 910 921
rect 1007 912 1012 917
rect 1114 912 1119 917
rect 1221 912 1226 917
rect 1328 912 1333 917
rect 1007 893 1012 898
rect 1114 893 1119 898
rect 1221 893 1226 898
rect 1328 893 1333 898
rect 447 800 452 805
rect -76 769 -71 774
rect 447 744 452 749
rect 437 737 442 742
rect 905 783 910 788
rect 1012 783 1017 788
rect 1119 783 1124 788
rect 1226 783 1231 788
rect 644 737 649 742
rect 905 740 910 745
rect 1007 736 1012 741
rect 1114 736 1119 741
rect 1221 736 1226 741
rect 1328 736 1333 741
rect 1007 717 1012 722
rect 1114 717 1119 722
rect 1221 717 1226 722
rect 1328 717 1333 722
rect 447 624 452 629
rect -76 593 -71 598
rect 447 568 452 573
rect 437 561 442 566
rect 905 607 910 612
rect 1012 607 1017 612
rect 1119 607 1124 612
rect 1226 607 1231 612
rect 644 561 649 566
rect 905 564 910 569
rect 1007 560 1012 565
rect 1114 560 1119 565
rect 1221 560 1226 565
rect 1328 560 1333 565
rect 1007 541 1012 546
rect 1114 541 1119 546
rect 1221 541 1226 546
rect 1328 541 1333 546
<< m4contact >>
rect 684 1856 689 1861
rect 165 1793 170 1798
rect 726 1805 731 1820
rect 206 1770 211 1775
rect 447 1770 452 1775
rect 1007 1815 1012 1820
rect 684 1773 689 1778
rect 684 1680 689 1685
rect 165 1617 170 1622
rect 726 1629 731 1644
rect 206 1594 211 1599
rect 447 1594 452 1599
rect 1007 1639 1012 1644
rect 684 1597 689 1602
rect 684 1504 689 1509
rect 165 1441 170 1446
rect 726 1453 731 1468
rect 206 1418 211 1423
rect 447 1418 452 1423
rect 1007 1463 1012 1468
rect 684 1421 689 1426
rect 684 1328 689 1333
rect 165 1265 170 1270
rect 726 1277 731 1292
rect 206 1242 211 1247
rect 447 1242 452 1247
rect 1007 1287 1012 1292
rect 684 1245 689 1250
rect 684 1152 689 1157
rect 165 1089 170 1094
rect 726 1101 731 1116
rect 206 1066 211 1071
rect 447 1066 452 1071
rect 1007 1111 1012 1116
rect 684 1069 689 1074
rect 684 976 689 981
rect 165 913 170 918
rect 726 925 731 940
rect 206 890 211 895
rect 447 890 452 895
rect 1007 935 1012 940
rect 684 893 689 898
rect 684 800 689 805
rect 165 737 170 742
rect 726 749 731 764
rect 206 714 211 719
rect 447 714 452 719
rect 1007 759 1012 764
rect 684 717 689 722
rect 684 624 689 629
rect 165 561 170 566
rect 726 573 731 588
rect 206 538 211 543
rect 447 538 452 543
rect 1007 583 1012 588
rect 684 541 689 546
<< metal4 >>
rect 452 1856 684 1861
rect 910 1839 1012 1844
rect 1017 1839 1119 1844
rect 1124 1839 1226 1844
rect 447 1805 726 1810
rect 731 1815 1007 1820
rect 170 1793 437 1798
rect 905 1793 910 1796
rect 437 1788 910 1793
rect 1012 1792 1114 1797
rect 1119 1792 1221 1797
rect 1226 1792 1328 1797
rect 211 1770 447 1775
rect 689 1773 1007 1778
rect 1012 1773 1114 1778
rect 1119 1773 1221 1778
rect 1226 1773 1328 1778
rect 452 1680 684 1685
rect 910 1663 1012 1668
rect 1017 1663 1119 1668
rect 1124 1663 1226 1668
rect 447 1629 726 1634
rect 731 1639 1007 1644
rect 170 1617 437 1622
rect 905 1617 910 1620
rect 437 1612 910 1617
rect 1012 1616 1114 1621
rect 1119 1616 1221 1621
rect 1226 1616 1328 1621
rect 211 1594 447 1599
rect 689 1597 1007 1602
rect 1012 1597 1114 1602
rect 1119 1597 1221 1602
rect 1226 1597 1328 1602
rect 452 1504 684 1509
rect 910 1487 1012 1492
rect 1017 1487 1119 1492
rect 1124 1487 1226 1492
rect 447 1453 726 1458
rect 731 1463 1007 1468
rect 170 1441 437 1446
rect 905 1441 910 1444
rect 437 1436 910 1441
rect 1012 1440 1114 1445
rect 1119 1440 1221 1445
rect 1226 1440 1328 1445
rect 211 1418 447 1423
rect 689 1421 1007 1426
rect 1012 1421 1114 1426
rect 1119 1421 1221 1426
rect 1226 1421 1328 1426
rect 452 1328 684 1333
rect 910 1311 1012 1316
rect 1017 1311 1119 1316
rect 1124 1311 1226 1316
rect 447 1277 726 1282
rect 731 1287 1007 1292
rect 170 1265 437 1270
rect 905 1265 910 1268
rect 437 1260 910 1265
rect 1012 1264 1114 1269
rect 1119 1264 1221 1269
rect 1226 1264 1328 1269
rect 211 1242 447 1247
rect 689 1245 1007 1250
rect 1012 1245 1114 1250
rect 1119 1245 1221 1250
rect 1226 1245 1328 1250
rect 452 1152 684 1157
rect 910 1135 1012 1140
rect 1017 1135 1119 1140
rect 1124 1135 1226 1140
rect 447 1101 726 1106
rect 731 1111 1007 1116
rect 170 1089 437 1094
rect 905 1089 910 1092
rect 437 1084 910 1089
rect 1012 1088 1114 1093
rect 1119 1088 1221 1093
rect 1226 1088 1328 1093
rect 211 1066 447 1071
rect 689 1069 1007 1074
rect 1012 1069 1114 1074
rect 1119 1069 1221 1074
rect 1226 1069 1328 1074
rect 452 976 684 981
rect 910 959 1012 964
rect 1017 959 1119 964
rect 1124 959 1226 964
rect 447 925 726 930
rect 731 935 1007 940
rect 170 913 437 918
rect 905 913 910 916
rect 437 908 910 913
rect 1012 912 1114 917
rect 1119 912 1221 917
rect 1226 912 1328 917
rect 211 890 447 895
rect 689 893 1007 898
rect 1012 893 1114 898
rect 1119 893 1221 898
rect 1226 893 1328 898
rect 452 800 684 805
rect 910 783 1012 788
rect 1017 783 1119 788
rect 1124 783 1226 788
rect 447 749 726 754
rect 731 759 1007 764
rect 170 737 437 742
rect 905 737 910 740
rect 437 732 910 737
rect 1012 736 1114 741
rect 1119 736 1221 741
rect 1226 736 1328 741
rect 211 714 447 719
rect 689 717 1007 722
rect 1012 717 1114 722
rect 1119 717 1221 722
rect 1226 717 1328 722
rect 452 624 684 629
rect 910 607 1012 612
rect 1017 607 1119 612
rect 1124 607 1226 612
rect 447 573 726 578
rect 731 583 1007 588
rect 170 561 437 566
rect 905 561 910 564
rect 437 556 910 561
rect 1012 560 1114 565
rect 1119 560 1221 565
rect 1226 560 1328 565
rect 211 538 447 543
rect 689 541 1007 546
rect 1012 541 1114 546
rect 1119 541 1221 546
rect 1226 541 1328 546
use latch  latch_4
timestamp 1765416915
transform -1 0 -351 0 1 463
box -392 82 -333 1369
use staticizer  staticizer_1
timestamp 1765334200
transform -1 0 43 0 1 1753
box 61 -1215 120 78
use latch  latch_0
timestamp 1765416915
transform 1 0 445 0 1 463
box -392 82 -333 1369
use staticizer  staticizer_0
timestamp 1765334200
transform 1 0 51 0 1 1753
box 61 -1215 120 78
use shift  shift_0
timestamp 1765416915
transform 1 0 330 0 1 2153
box -138 -1615 46 -268
use latch  latch_3
timestamp 1765416915
transform 1 0 768 0 1 456
box -392 82 -333 1369
use fblock  fblock_0
timestamp 1765416915
transform 1 0 535 0 1 2993
box -80 -2455 50 -1047
use addsub  addsub_0
timestamp 1765338694
transform 1 0 675 0 1 712
box -14 -174 166 1225
use latch  latch_1
timestamp 1765416915
transform 1 0 975 0 1 456
box -392 82 -333 1369
use latch  latch_2
timestamp 1765416915
transform 1 0 1236 0 1 459
box -392 82 -333 1369
use reg  reg_0
timestamp 1765316199
transform 1 0 928 0 1 936
box -14 -398 76 940
use reg  reg_1
timestamp 1765316199
transform 1 0 1035 0 1 936
box -14 -398 76 940
use reg  reg_2
timestamp 1765316199
transform 1 0 1142 0 1 936
box -14 -398 76 940
use reg  reg_3
timestamp 1765316199
transform 1 0 1249 0 1 936
box -14 -398 76 940
<< end >>
