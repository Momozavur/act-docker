magic
tech scmos
timestamp 1765745113
<< polysilicon >>
rect 924 2012 946 2014
rect 921 1939 923 1989
rect 148 1893 159 1895
rect 835 1893 842 1895
rect 1710 1893 1716 1895
rect 2510 1893 2516 1895
rect 148 1883 159 1885
rect 148 1873 159 1875
rect 1619 1865 1621 1867
rect 96 1840 98 1862
rect 37 1805 38 1808
rect 1550 1808 1553 1813
rect 52 1805 53 1808
rect 678 1804 679 1806
rect 37 1629 38 1632
rect 1550 1632 1553 1637
rect 52 1629 53 1632
rect 678 1628 679 1630
rect 37 1453 38 1456
rect 1550 1456 1553 1461
rect 52 1453 53 1456
rect 678 1452 679 1454
rect 37 1277 38 1280
rect 1550 1280 1553 1285
rect 52 1277 53 1280
rect 678 1276 679 1278
rect 37 1101 38 1104
rect 1550 1104 1553 1109
rect 52 1101 53 1104
rect 678 1100 679 1102
rect 37 925 38 928
rect 1550 928 1553 933
rect 52 925 53 928
rect 678 924 679 926
rect 37 749 38 752
rect 1550 752 1553 757
rect 52 749 53 752
rect 678 748 679 750
rect 37 573 38 576
rect 1550 576 1553 581
rect 52 573 53 576
rect 678 572 679 574
<< polycontact >>
rect 919 2009 924 2014
rect 860 1991 865 1996
rect 918 1989 923 1994
rect 957 1989 962 1994
rect 857 1939 862 1944
rect 919 1934 924 1939
rect 842 1893 847 1898
rect 1606 1874 1611 1879
rect 2406 1874 2411 1879
rect 96 1835 101 1840
rect 1545 1808 1550 1813
rect -24 1800 -19 1805
rect 109 1800 114 1805
rect 1776 1804 1781 1809
rect 2351 1801 2356 1806
rect 2575 1804 2580 1809
rect 2699 1804 2704 1809
rect 2823 1804 2828 1809
rect 373 1796 378 1801
rect 580 1795 585 1800
rect 2640 1799 2645 1804
rect 2764 1799 2769 1804
rect 1606 1698 1611 1703
rect 2406 1698 2411 1703
rect 1545 1632 1550 1637
rect -24 1624 -19 1629
rect 109 1624 114 1629
rect 1776 1628 1781 1633
rect 2351 1625 2356 1630
rect 2575 1628 2580 1633
rect 2699 1628 2704 1633
rect 2823 1628 2828 1633
rect 373 1620 378 1625
rect 580 1619 585 1624
rect 2640 1623 2645 1628
rect 2764 1623 2769 1628
rect 1606 1522 1611 1527
rect 2406 1522 2411 1527
rect 1545 1456 1550 1461
rect -24 1448 -19 1453
rect 109 1448 114 1453
rect 1776 1452 1781 1457
rect 2351 1449 2356 1454
rect 2575 1452 2580 1457
rect 2699 1452 2704 1457
rect 2823 1452 2828 1457
rect 373 1444 378 1449
rect 580 1443 585 1448
rect 2640 1447 2645 1452
rect 2764 1447 2769 1452
rect 1606 1346 1611 1351
rect 2406 1346 2411 1351
rect 1545 1280 1550 1285
rect -24 1272 -19 1277
rect 109 1272 114 1277
rect 1776 1276 1781 1281
rect 2351 1273 2356 1278
rect 2575 1276 2580 1281
rect 2699 1276 2704 1281
rect 2823 1276 2828 1281
rect 373 1268 378 1273
rect 580 1267 585 1272
rect 2640 1271 2645 1276
rect 2764 1271 2769 1276
rect 1606 1170 1611 1175
rect 2406 1170 2411 1175
rect 1545 1104 1550 1109
rect -24 1096 -19 1101
rect 109 1096 114 1101
rect 1776 1100 1781 1105
rect 2351 1097 2356 1102
rect 2575 1100 2580 1105
rect 2699 1100 2704 1105
rect 2823 1100 2828 1105
rect 373 1092 378 1097
rect 580 1091 585 1096
rect 2640 1095 2645 1100
rect 2764 1095 2769 1100
rect 1606 994 1611 999
rect 2406 994 2411 999
rect 1545 928 1550 933
rect -24 920 -19 925
rect 109 920 114 925
rect 1776 924 1781 929
rect 2351 921 2356 926
rect 2575 924 2580 929
rect 2699 924 2704 929
rect 2823 924 2828 929
rect 373 916 378 921
rect 580 915 585 920
rect 2640 919 2645 924
rect 2764 919 2769 924
rect 1606 818 1611 823
rect 2406 818 2411 823
rect 1545 752 1550 757
rect -24 744 -19 749
rect 109 744 114 749
rect 1776 748 1781 753
rect 2351 745 2356 750
rect 2575 748 2580 753
rect 2699 748 2704 753
rect 2823 748 2828 753
rect 373 740 378 745
rect 580 739 585 744
rect 2640 743 2645 748
rect 2764 743 2769 748
rect 1606 642 1611 647
rect 2406 642 2411 647
rect 1545 576 1550 581
rect -24 568 -19 573
rect 109 568 114 573
rect 1776 572 1781 577
rect 2351 569 2356 574
rect 2575 572 2580 577
rect 2699 572 2704 577
rect 2823 572 2828 577
rect 373 564 378 569
rect 580 563 585 568
rect 2640 567 2645 572
rect 2764 567 2769 572
<< metal1 >>
rect 860 1969 865 1991
rect 1404 1990 1409 1996
rect 1904 1990 1909 1996
rect 2204 1991 2209 1996
rect 979 1961 984 1978
rect 985 1902 992 1907
rect 1380 1902 1385 1972
rect 842 1898 847 1901
rect 1422 1899 1427 1969
rect 1880 1902 1885 1972
rect 1922 1899 1927 1969
rect 2180 1902 2185 1972
rect 2222 1899 2227 1969
rect 1380 1876 1386 1882
rect 1422 1870 1427 1879
rect 1880 1876 1886 1882
rect 1796 1867 1807 1872
rect 1922 1870 1927 1879
rect 2180 1876 2186 1882
rect 2222 1870 2227 1879
rect 2596 1867 2607 1872
rect 2720 1867 2731 1872
rect 2844 1867 2855 1872
rect -51 1860 -33 1865
rect 65 1845 73 1851
rect 101 1835 105 1840
rect 136 1836 141 1856
rect 910 1844 915 1849
rect 1017 1844 1022 1849
rect 1124 1844 1129 1849
rect 1231 1844 1236 1849
rect -80 1825 -75 1830
rect 661 1829 666 1834
rect 1438 1825 1443 1846
rect 1536 1834 1546 1839
rect 1938 1825 1943 1846
rect 2037 1844 2042 1849
rect 2238 1825 2243 1846
rect 2336 1834 2350 1839
rect 1431 1820 1443 1825
rect 1931 1820 1943 1825
rect 2231 1820 2243 1825
rect 369 1796 373 1801
rect 369 1775 374 1796
rect 563 1795 580 1800
rect 1004 1787 1007 1792
rect 1111 1787 1114 1792
rect 1218 1787 1221 1792
rect 1325 1787 1328 1792
rect 1431 1779 1436 1820
rect 1776 1796 1781 1804
rect 1525 1787 1527 1792
rect 1931 1779 1936 1820
rect 2025 1787 2028 1792
rect 2132 1787 2135 1792
rect 2231 1779 2236 1820
rect 2575 1796 2580 1804
rect 2699 1796 2704 1804
rect 2823 1796 2828 1804
rect 2325 1787 2328 1792
rect 363 1770 374 1775
rect 1409 1774 1436 1779
rect 1909 1774 1936 1779
rect 2209 1774 2236 1779
rect 1551 1741 1556 1760
rect 910 1668 915 1673
rect 1017 1668 1022 1673
rect 1124 1668 1129 1673
rect 1231 1668 1236 1673
rect -80 1649 -75 1654
rect 1438 1649 1443 1670
rect 1938 1649 1943 1670
rect 2037 1668 2042 1673
rect 2238 1649 2243 1670
rect 1431 1644 1443 1649
rect 1931 1644 1943 1649
rect 2231 1644 2243 1649
rect 369 1620 373 1625
rect 369 1599 374 1620
rect 563 1619 580 1624
rect 1004 1611 1007 1616
rect 1111 1611 1114 1616
rect 1218 1611 1221 1616
rect 1325 1611 1328 1616
rect 1431 1603 1436 1644
rect 1776 1620 1781 1628
rect 1525 1611 1527 1616
rect 1931 1603 1936 1644
rect 2025 1611 2028 1616
rect 2132 1611 2135 1616
rect 2231 1603 2236 1644
rect 2575 1620 2580 1628
rect 2699 1620 2704 1628
rect 2823 1620 2828 1628
rect 2325 1611 2328 1616
rect 363 1594 374 1599
rect 1409 1598 1436 1603
rect 1909 1598 1936 1603
rect 2209 1598 2236 1603
rect 910 1492 915 1497
rect 1017 1492 1022 1497
rect 1124 1492 1129 1497
rect 1231 1492 1236 1497
rect -80 1473 -75 1478
rect 1438 1473 1443 1494
rect 1938 1473 1943 1494
rect 2037 1492 2042 1497
rect 2238 1473 2243 1494
rect 1431 1468 1443 1473
rect 1931 1468 1943 1473
rect 2231 1468 2243 1473
rect 369 1444 373 1449
rect 369 1423 374 1444
rect 563 1443 580 1448
rect 1004 1435 1007 1440
rect 1111 1435 1114 1440
rect 1218 1435 1221 1440
rect 1325 1435 1328 1440
rect 1431 1427 1436 1468
rect 1776 1444 1781 1452
rect 1525 1435 1527 1440
rect 1931 1427 1936 1468
rect 2025 1435 2028 1440
rect 2132 1435 2135 1440
rect 2231 1427 2236 1468
rect 2575 1444 2580 1452
rect 2699 1444 2704 1452
rect 2823 1444 2828 1452
rect 2325 1435 2328 1440
rect 363 1418 374 1423
rect 1409 1422 1436 1427
rect 1909 1422 1936 1427
rect 2209 1422 2236 1427
rect 910 1316 915 1321
rect 1017 1316 1022 1321
rect 1124 1316 1129 1321
rect 1231 1316 1236 1321
rect -80 1297 -75 1302
rect 1438 1297 1443 1318
rect 1938 1297 1943 1318
rect 2037 1316 2042 1321
rect 2238 1297 2243 1318
rect 1431 1292 1443 1297
rect 1931 1292 1943 1297
rect 2231 1292 2243 1297
rect 369 1268 373 1273
rect 369 1247 374 1268
rect 563 1267 580 1272
rect 1004 1259 1007 1264
rect 1111 1259 1114 1264
rect 1218 1259 1221 1264
rect 1325 1259 1328 1264
rect 1431 1251 1436 1292
rect 1776 1268 1781 1276
rect 1525 1259 1527 1264
rect 1931 1251 1936 1292
rect 2025 1259 2028 1264
rect 2132 1259 2135 1264
rect 2231 1251 2236 1292
rect 2575 1268 2580 1276
rect 2699 1268 2704 1276
rect 2823 1268 2828 1276
rect 2325 1259 2328 1264
rect 363 1242 374 1247
rect 1409 1246 1436 1251
rect 1909 1246 1936 1251
rect 2209 1246 2236 1251
rect 910 1140 915 1145
rect 1017 1140 1022 1145
rect 1124 1140 1129 1145
rect 1231 1140 1236 1145
rect -80 1121 -75 1126
rect 1438 1121 1443 1142
rect 1938 1121 1943 1142
rect 2037 1140 2042 1145
rect 2238 1121 2243 1142
rect 1431 1116 1443 1121
rect 1931 1116 1943 1121
rect 2231 1116 2243 1121
rect 369 1092 373 1097
rect 369 1071 374 1092
rect 563 1091 580 1096
rect 1004 1083 1007 1088
rect 1111 1083 1114 1088
rect 1218 1083 1221 1088
rect 1325 1083 1328 1088
rect 1431 1075 1436 1116
rect 1776 1092 1781 1100
rect 1525 1083 1527 1088
rect 1931 1075 1936 1116
rect 2025 1083 2028 1088
rect 2132 1083 2135 1088
rect 2231 1075 2236 1116
rect 2575 1092 2580 1100
rect 2699 1092 2704 1100
rect 2823 1092 2828 1100
rect 2325 1083 2328 1088
rect 363 1066 374 1071
rect 1409 1070 1436 1075
rect 1909 1070 1936 1075
rect 2209 1070 2236 1075
rect 910 964 915 969
rect 1017 964 1022 969
rect 1124 964 1129 969
rect 1231 964 1236 969
rect -80 945 -75 950
rect 1438 945 1443 966
rect 1938 945 1943 966
rect 2037 964 2042 969
rect 2238 945 2243 966
rect 1431 940 1443 945
rect 1931 940 1943 945
rect 2231 940 2243 945
rect 369 916 373 921
rect 369 895 374 916
rect 563 915 580 920
rect 1004 907 1007 912
rect 1111 907 1114 912
rect 1218 907 1221 912
rect 1325 907 1328 912
rect 1431 899 1436 940
rect 1776 916 1781 924
rect 1525 907 1527 912
rect 1931 899 1936 940
rect 2025 907 2028 912
rect 2132 907 2135 912
rect 2231 899 2236 940
rect 2575 916 2580 924
rect 2699 916 2704 924
rect 2823 916 2828 924
rect 2325 907 2328 912
rect 363 890 374 895
rect 1409 894 1436 899
rect 1909 894 1936 899
rect 2209 894 2236 899
rect 910 788 915 793
rect 1017 788 1022 793
rect 1124 788 1129 793
rect 1231 788 1236 793
rect -80 769 -75 774
rect 1438 769 1443 790
rect 1938 769 1943 790
rect 2037 788 2042 793
rect 2238 769 2243 790
rect 1431 764 1443 769
rect 1931 764 1943 769
rect 2231 764 2243 769
rect 369 740 373 745
rect 369 719 374 740
rect 563 739 580 744
rect 1004 731 1007 736
rect 1111 731 1114 736
rect 1218 731 1221 736
rect 1325 731 1328 736
rect 1431 723 1436 764
rect 1776 740 1781 748
rect 1525 731 1527 736
rect 1931 723 1936 764
rect 2025 731 2028 736
rect 2132 731 2135 736
rect 2231 723 2236 764
rect 2575 740 2580 748
rect 2699 740 2704 748
rect 2823 740 2828 748
rect 2325 731 2328 736
rect 363 714 374 719
rect 1409 718 1436 723
rect 1909 718 1936 723
rect 2209 718 2236 723
rect 910 612 915 617
rect 1017 612 1022 617
rect 1124 612 1129 617
rect 1231 612 1236 617
rect -80 593 -75 598
rect 1438 593 1443 614
rect 1938 593 1943 614
rect 2037 612 2042 617
rect 2238 593 2243 614
rect 1431 588 1443 593
rect 1931 588 1943 593
rect 2231 588 2243 593
rect 369 564 373 569
rect 369 543 374 564
rect 563 563 580 568
rect 1004 555 1007 560
rect 1111 555 1114 560
rect 1218 555 1221 560
rect 1325 555 1328 560
rect 1431 547 1436 588
rect 1776 564 1781 572
rect 1525 555 1527 560
rect 1931 547 1936 588
rect 2025 555 2028 560
rect 2132 555 2135 560
rect 2231 547 2236 588
rect 2345 569 2351 581
rect 2575 564 2580 572
rect 2699 564 2704 572
rect 2823 564 2828 572
rect 2325 555 2328 560
rect 363 538 374 543
rect 1409 542 1436 547
rect 1909 542 1936 547
rect 2209 542 2236 547
<< m2contact >>
rect 927 2013 932 2018
rect 924 1954 929 1959
rect 1623 1916 1628 1921
rect 452 1856 457 1861
rect 1343 1850 1348 1855
rect 1843 1850 1848 1855
rect 2143 1850 2148 1855
rect 905 1844 910 1849
rect 1012 1844 1017 1849
rect 1119 1844 1124 1849
rect 1226 1844 1231 1849
rect 2032 1844 2037 1849
rect 432 1793 437 1798
rect 452 1795 457 1800
rect 639 1793 644 1798
rect 900 1796 905 1801
rect 1007 1787 1012 1792
rect 1114 1787 1119 1792
rect 1221 1787 1226 1792
rect 1328 1787 1333 1792
rect 1343 1791 1348 1796
rect 1527 1787 1532 1792
rect 1849 1791 1854 1796
rect 2028 1787 2033 1792
rect 2143 1791 2148 1796
rect 2626 1801 2631 1806
rect 2328 1787 2333 1792
rect 833 1741 838 1762
rect 1546 1741 1551 1760
rect 2346 1741 2351 1760
rect 739 1711 744 1732
rect 1614 1711 1619 1732
rect 2414 1711 2419 1732
rect 452 1680 457 1685
rect 1343 1674 1348 1679
rect 1843 1674 1848 1679
rect 2143 1674 2148 1679
rect 905 1668 910 1673
rect 1012 1668 1017 1673
rect 1119 1668 1124 1673
rect 1226 1668 1231 1673
rect 2032 1668 2037 1673
rect 432 1617 437 1622
rect 452 1619 457 1624
rect 639 1617 644 1622
rect 900 1620 905 1625
rect 1007 1611 1012 1616
rect 1114 1611 1119 1616
rect 1221 1611 1226 1616
rect 1328 1611 1333 1616
rect 1343 1615 1348 1620
rect 1527 1611 1532 1616
rect 1849 1615 1854 1620
rect 2028 1611 2033 1616
rect 2143 1615 2148 1620
rect 2626 1625 2631 1630
rect 2328 1611 2333 1616
rect 452 1504 457 1509
rect 1343 1498 1348 1503
rect 1843 1498 1848 1503
rect 2143 1498 2148 1503
rect 905 1492 910 1497
rect 1012 1492 1017 1497
rect 1119 1492 1124 1497
rect 1226 1492 1231 1497
rect 2032 1492 2037 1497
rect 432 1441 437 1446
rect 452 1443 457 1448
rect 639 1441 644 1446
rect 900 1444 905 1449
rect 1007 1435 1012 1440
rect 1114 1435 1119 1440
rect 1221 1435 1226 1440
rect 1328 1435 1333 1440
rect 1343 1439 1348 1444
rect 1527 1435 1532 1440
rect 1849 1439 1854 1444
rect 2028 1435 2033 1440
rect 2143 1439 2148 1444
rect 2626 1449 2631 1454
rect 2328 1435 2333 1440
rect 452 1328 457 1333
rect 1343 1322 1348 1327
rect 1843 1322 1848 1327
rect 2143 1322 2148 1327
rect 905 1316 910 1321
rect 1012 1316 1017 1321
rect 1119 1316 1124 1321
rect 1226 1316 1231 1321
rect 2032 1316 2037 1321
rect 432 1265 437 1270
rect 452 1267 457 1272
rect 639 1265 644 1270
rect 900 1268 905 1273
rect 1007 1259 1012 1264
rect 1114 1259 1119 1264
rect 1221 1259 1226 1264
rect 1328 1259 1333 1264
rect 1343 1263 1348 1268
rect 1527 1259 1532 1264
rect 1849 1263 1854 1268
rect 2028 1259 2033 1264
rect 2143 1263 2148 1268
rect 2626 1273 2631 1278
rect 2328 1259 2333 1264
rect 452 1152 457 1157
rect 1343 1146 1348 1151
rect 1843 1146 1848 1151
rect 2143 1146 2148 1151
rect 905 1140 910 1145
rect 1012 1140 1017 1145
rect 1119 1140 1124 1145
rect 1226 1140 1231 1145
rect 2032 1140 2037 1145
rect 432 1089 437 1094
rect 452 1091 457 1096
rect 639 1089 644 1094
rect 900 1092 905 1097
rect 1007 1083 1012 1088
rect 1114 1083 1119 1088
rect 1221 1083 1226 1088
rect 1328 1083 1333 1088
rect 1343 1087 1348 1092
rect 1527 1083 1532 1088
rect 1849 1087 1854 1092
rect 2028 1083 2033 1088
rect 2143 1087 2148 1092
rect 2626 1097 2631 1102
rect 2328 1083 2333 1088
rect 452 976 457 981
rect 1343 970 1348 975
rect 1843 970 1848 975
rect 2143 970 2148 975
rect 905 964 910 969
rect 1012 964 1017 969
rect 1119 964 1124 969
rect 1226 964 1231 969
rect 2032 964 2037 969
rect 432 913 437 918
rect 452 915 457 920
rect 639 913 644 918
rect 900 916 905 921
rect 1007 907 1012 912
rect 1114 907 1119 912
rect 1221 907 1226 912
rect 1328 907 1333 912
rect 1343 911 1348 916
rect 1527 907 1532 912
rect 1849 911 1854 916
rect 2028 907 2033 912
rect 2143 911 2148 916
rect 2626 921 2631 926
rect 2328 907 2333 912
rect 452 800 457 805
rect 1343 794 1348 799
rect 1843 794 1848 799
rect 2143 794 2148 799
rect 905 788 910 793
rect 1012 788 1017 793
rect 1119 788 1124 793
rect 1226 788 1231 793
rect 2032 788 2037 793
rect 432 737 437 742
rect 452 739 457 744
rect 639 737 644 742
rect 900 740 905 745
rect 1007 731 1012 736
rect 1114 731 1119 736
rect 1221 731 1226 736
rect 1328 731 1333 736
rect 1343 735 1348 740
rect 1527 731 1532 736
rect 1849 735 1854 740
rect 2028 731 2033 736
rect 2143 735 2148 740
rect 2626 745 2631 750
rect 2328 731 2333 736
rect 452 624 457 629
rect 1343 618 1348 623
rect 1843 618 1848 623
rect 2143 618 2148 623
rect 905 612 910 617
rect 1012 612 1017 617
rect 1119 612 1124 617
rect 1226 612 1231 617
rect 2032 612 2037 617
rect 432 561 437 566
rect 452 563 457 568
rect 639 561 644 566
rect 900 564 905 569
rect 1007 555 1012 560
rect 1114 555 1119 560
rect 1221 555 1226 560
rect 1328 555 1333 560
rect 1343 559 1348 564
rect 1527 555 1532 560
rect 1849 559 1854 564
rect 2028 555 2033 560
rect 2143 559 2148 564
rect 2626 569 2631 574
rect 2328 555 2333 560
<< pm12contact >>
rect 159 1893 164 1898
rect 1716 1893 1721 1898
rect 2516 1893 2521 1898
rect 159 1882 164 1887
rect 159 1870 164 1875
rect 731 1874 736 1879
rect 38 1805 43 1810
rect 47 1805 52 1810
rect 679 1801 684 1806
rect 841 1801 846 1806
rect 1716 1801 1721 1806
rect 2516 1801 2521 1806
rect 731 1698 736 1703
rect 38 1629 43 1634
rect 47 1629 52 1634
rect 679 1625 684 1630
rect 841 1625 846 1630
rect 1716 1625 1721 1630
rect 2516 1625 2521 1630
rect 731 1522 736 1527
rect 38 1453 43 1458
rect 47 1453 52 1458
rect 679 1449 684 1454
rect 841 1449 846 1454
rect 1716 1449 1721 1454
rect 2516 1449 2521 1454
rect 731 1346 736 1351
rect 38 1277 43 1282
rect 47 1277 52 1282
rect 679 1273 684 1278
rect 841 1273 846 1278
rect 1716 1273 1721 1278
rect 2516 1273 2521 1278
rect 731 1170 736 1175
rect 38 1101 43 1106
rect 47 1101 52 1106
rect 679 1097 684 1102
rect 841 1097 846 1102
rect 1716 1097 1721 1102
rect 2516 1097 2521 1102
rect 731 994 736 999
rect 38 925 43 930
rect 47 925 52 930
rect 679 921 684 926
rect 841 921 846 926
rect 1716 921 1721 926
rect 2516 921 2521 926
rect 731 818 736 823
rect 38 749 43 754
rect 47 749 52 754
rect 679 745 684 750
rect 841 745 846 750
rect 1716 745 1721 750
rect 2516 745 2521 750
rect 731 642 736 647
rect 38 573 43 578
rect 47 573 52 578
rect 679 569 684 574
rect 841 569 846 574
rect 1716 569 1721 574
rect 2516 569 2521 574
<< metal2 >>
rect 870 2013 927 2018
rect 870 1959 1000 1962
rect 870 1958 924 1959
rect 865 1957 924 1958
rect 929 1957 1000 1959
rect 986 1941 991 1957
rect 1628 1916 1721 1921
rect 957 1914 1004 1916
rect 952 1911 1004 1914
rect 980 1900 985 1905
rect 1058 1902 1063 1907
rect 1716 1898 1721 1916
rect 914 1876 919 1880
rect 1021 1876 1026 1880
rect 1128 1876 1133 1880
rect 1235 1876 1240 1880
rect 1435 1876 1440 1879
rect 1935 1876 1940 1879
rect 2042 1876 2047 1880
rect 2235 1876 2240 1880
rect 1492 1844 1496 1849
rect 1704 1801 1708 1806
rect 447 1795 452 1800
rect 1532 1787 1601 1792
rect 2333 1787 2401 1792
rect 1002 1773 1007 1778
rect 1109 1773 1114 1778
rect 1216 1773 1221 1778
rect 1323 1773 1328 1778
rect 1523 1773 1528 1778
rect 2023 1773 2033 1778
rect 2130 1773 2135 1778
rect 2323 1773 2333 1778
rect 2028 1769 2033 1773
rect 2328 1769 2333 1773
rect 1492 1668 1496 1673
rect 1704 1625 1708 1630
rect 447 1619 452 1624
rect 1532 1611 1601 1616
rect 2333 1611 2401 1616
rect 1002 1597 1007 1602
rect 1109 1597 1114 1602
rect 1216 1597 1221 1602
rect 1323 1597 1328 1602
rect 1523 1597 1528 1602
rect 2023 1597 2033 1602
rect 2130 1597 2135 1602
rect 2323 1597 2333 1602
rect 2028 1593 2033 1597
rect 2328 1593 2333 1597
rect 1492 1492 1496 1497
rect 1704 1449 1708 1454
rect 447 1443 452 1448
rect 1532 1435 1601 1440
rect 2333 1435 2401 1440
rect 1002 1421 1007 1426
rect 1109 1421 1114 1426
rect 1216 1421 1221 1426
rect 1323 1421 1328 1426
rect 1523 1421 1528 1426
rect 2023 1421 2033 1426
rect 2130 1421 2135 1426
rect 2323 1421 2333 1426
rect 2028 1417 2033 1421
rect 2328 1417 2333 1421
rect 1492 1316 1496 1321
rect 1704 1273 1708 1278
rect 447 1267 452 1272
rect 1532 1259 1601 1264
rect 2333 1259 2401 1264
rect 1002 1245 1007 1250
rect 1109 1245 1114 1250
rect 1216 1245 1221 1250
rect 1323 1245 1328 1250
rect 1523 1245 1528 1250
rect 2023 1245 2033 1250
rect 2130 1245 2135 1250
rect 2323 1245 2333 1250
rect 2028 1241 2033 1245
rect 2328 1241 2333 1245
rect 1492 1140 1496 1145
rect 1704 1097 1708 1102
rect 447 1091 452 1096
rect 1532 1083 1601 1088
rect 2333 1083 2401 1088
rect 1002 1069 1007 1074
rect 1109 1069 1114 1074
rect 1216 1069 1221 1074
rect 1323 1069 1328 1074
rect 1523 1069 1528 1074
rect 2023 1069 2033 1074
rect 2130 1069 2135 1074
rect 2323 1069 2333 1074
rect 2028 1065 2033 1069
rect 2328 1065 2333 1069
rect 1492 964 1496 969
rect 1704 921 1708 926
rect 447 915 452 920
rect 1532 907 1601 912
rect 2333 907 2401 912
rect 1002 893 1007 898
rect 1109 893 1114 898
rect 1216 893 1221 898
rect 1323 893 1328 898
rect 1523 893 1528 898
rect 2023 893 2033 898
rect 2130 893 2135 898
rect 2323 893 2333 898
rect 2028 889 2033 893
rect 2328 889 2333 893
rect 1492 788 1496 793
rect 1704 745 1708 750
rect 447 739 452 744
rect 1532 731 1601 736
rect 2333 731 2401 736
rect 1002 717 1007 722
rect 1109 717 1114 722
rect 1216 717 1221 722
rect 1323 717 1328 722
rect 1523 717 1528 722
rect 2023 717 2033 722
rect 2130 717 2135 722
rect 2323 717 2333 722
rect 2028 713 2033 717
rect 2328 713 2333 717
rect 1492 612 1496 617
rect 836 569 841 574
rect 1704 569 1708 574
rect 1711 569 1716 574
rect 2511 569 2516 574
rect 447 563 452 568
rect 1532 555 1601 560
rect 2333 555 2401 560
rect 1002 541 1007 546
rect 1109 541 1114 546
rect 1216 541 1221 546
rect 1323 541 1328 546
rect 1523 541 1528 546
rect 2023 541 2033 546
rect 2130 541 2135 546
rect 2323 541 2333 546
rect 2028 537 2033 541
rect 2328 537 2333 541
<< m3contact >>
rect 726 1874 731 1879
rect 38 1800 43 1805
rect 684 1801 689 1806
rect 1601 1787 1606 1792
rect 2401 1787 2406 1792
rect 726 1698 731 1703
rect 38 1624 43 1629
rect 684 1625 689 1630
rect 1601 1611 1606 1616
rect 2401 1611 2406 1616
rect 726 1522 731 1527
rect 38 1448 43 1453
rect 684 1449 689 1454
rect 1601 1435 1606 1440
rect 2401 1435 2406 1440
rect 726 1346 731 1351
rect 38 1272 43 1277
rect 684 1273 689 1278
rect 1601 1259 1606 1264
rect 2401 1259 2406 1264
rect 726 1170 731 1175
rect 38 1096 43 1101
rect 684 1097 689 1102
rect 1601 1083 1606 1088
rect 2401 1083 2406 1088
rect 726 994 731 999
rect 38 920 43 925
rect 684 921 689 926
rect 1601 907 1606 912
rect 2401 907 2406 912
rect 726 818 731 823
rect 38 744 43 749
rect 684 745 689 750
rect 1601 731 1606 736
rect 2401 731 2406 736
rect 726 642 731 647
rect 38 568 43 573
rect 684 569 689 574
rect 1601 555 1606 560
rect 2401 555 2406 560
<< m123contact >>
rect 865 2013 870 2018
rect 919 2004 924 2009
rect 962 1989 967 1994
rect 953 1971 958 1976
rect 877 1966 882 1971
rect 865 1958 870 1963
rect 852 1939 857 1944
rect 952 1914 957 1919
rect -30 1884 -25 1889
rect 1793 1885 1798 1890
rect 2593 1885 2598 1890
rect 2717 1885 2722 1890
rect 2841 1885 2846 1890
rect 1601 1874 1606 1879
rect 2401 1874 2406 1879
rect 1771 1867 1776 1872
rect 1807 1867 1812 1872
rect 2571 1867 2576 1872
rect 2607 1867 2612 1872
rect 2695 1867 2700 1872
rect 2731 1867 2736 1872
rect 2819 1867 2824 1872
rect 2855 1867 2860 1872
rect -56 1860 -51 1865
rect -20 1860 -15 1865
rect -42 1842 -37 1847
rect 150 1845 155 1850
rect 68 1840 73 1845
rect 105 1835 110 1840
rect 141 1836 146 1841
rect 1780 1843 1785 1848
rect 2580 1843 2585 1848
rect 2704 1843 2709 1848
rect 2828 1843 2833 1848
rect 160 1825 165 1830
rect 1820 1828 1825 1833
rect 2635 1799 2640 1804
rect 2759 1799 2764 1804
rect 1601 1698 1606 1703
rect 2401 1698 2406 1703
rect 160 1649 165 1654
rect 1820 1652 1825 1657
rect 2635 1623 2640 1628
rect 2759 1623 2764 1628
rect 1601 1522 1606 1527
rect 2401 1522 2406 1527
rect 160 1473 165 1478
rect 1820 1476 1825 1481
rect 2635 1447 2640 1452
rect 2759 1447 2764 1452
rect 1601 1346 1606 1351
rect 2401 1346 2406 1351
rect 160 1297 165 1302
rect 1820 1300 1825 1305
rect 2635 1271 2640 1276
rect 2759 1271 2764 1276
rect 1601 1170 1606 1175
rect 2401 1170 2406 1175
rect 160 1121 165 1126
rect 1820 1124 1825 1129
rect 2635 1095 2640 1100
rect 2759 1095 2764 1100
rect 1601 994 1606 999
rect 2401 994 2406 999
rect 160 945 165 950
rect 1820 948 1825 953
rect 2635 919 2640 924
rect 2759 919 2764 924
rect 1601 818 1606 823
rect 2401 818 2406 823
rect 160 769 165 774
rect 1820 772 1825 777
rect 2635 743 2640 748
rect 2759 743 2764 748
rect 1601 642 1606 647
rect 2401 642 2406 647
rect 160 593 165 598
rect 1820 596 1825 601
rect 2635 567 2640 572
rect 2759 567 2764 572
rect 812 538 817 543
rect 1687 537 1692 542
<< metal3 >>
rect 456 1922 461 1948
rect 488 1922 493 1948
rect 522 1922 527 1948
rect 555 1922 560 1948
rect -56 1831 -51 1860
rect -42 1831 -37 1842
rect -30 1831 -25 1884
rect 284 1885 289 1890
rect 346 1885 351 1890
rect 635 1887 640 1972
rect 865 1963 870 2013
rect 914 1977 919 2009
rect 1059 2000 1064 2005
rect 952 1971 953 1976
rect 870 1958 872 1963
rect -20 1831 -15 1860
rect 115 1845 150 1850
rect 68 1831 73 1840
rect 105 1831 110 1835
rect 115 1831 120 1845
rect 141 1831 146 1836
rect 38 1775 43 1800
rect 165 1798 170 1830
rect 428 1824 433 1870
rect 635 1824 640 1882
rect 812 1939 852 1944
rect 684 1806 689 1856
rect 447 1775 452 1800
rect 726 1820 731 1874
rect 684 1778 689 1801
rect 38 1599 43 1624
rect 165 1622 170 1654
rect 684 1630 689 1680
rect 447 1599 452 1624
rect 726 1644 731 1698
rect 684 1602 689 1625
rect 38 1423 43 1448
rect 165 1446 170 1478
rect 684 1454 689 1504
rect 447 1423 452 1448
rect 726 1468 731 1522
rect 684 1426 689 1449
rect 38 1247 43 1272
rect 165 1270 170 1302
rect 684 1278 689 1328
rect 447 1247 452 1272
rect 726 1292 731 1346
rect 684 1250 689 1273
rect 38 1071 43 1096
rect 165 1094 170 1126
rect 684 1102 689 1152
rect 447 1071 452 1096
rect 726 1116 731 1170
rect 684 1074 689 1097
rect 38 895 43 920
rect 165 918 170 950
rect 684 926 689 976
rect 447 895 452 920
rect 726 940 731 994
rect 684 898 689 921
rect 38 719 43 744
rect 165 742 170 774
rect 684 750 689 800
rect 447 719 452 744
rect 726 764 731 818
rect 684 722 689 745
rect 38 543 43 568
rect 165 566 170 598
rect 684 574 689 624
rect 447 543 452 568
rect 726 588 731 642
rect 684 546 689 569
rect 812 543 817 1939
rect 867 1889 872 1958
rect 847 1884 872 1889
rect 847 1827 852 1884
rect 877 1847 882 1966
rect 914 1917 919 1956
rect 859 1842 882 1847
rect 896 1912 919 1917
rect 952 1919 957 1971
rect 962 1961 967 1989
rect 896 1898 901 1912
rect 896 1868 901 1893
rect 925 1876 930 1880
rect 952 1876 957 1914
rect 998 1876 1003 1880
rect 1032 1876 1037 1880
rect 1105 1876 1110 1880
rect 1139 1876 1144 1880
rect 1212 1876 1217 1880
rect 1246 1876 1251 1880
rect 1319 1876 1324 1880
rect 1446 1876 1451 1879
rect 1519 1876 1524 1879
rect 859 1827 864 1842
rect 896 1827 901 1863
rect 905 1801 910 1839
rect 1007 1797 1012 1815
rect 1601 1792 1606 1874
rect 905 1625 910 1663
rect 1007 1621 1012 1639
rect 1601 1616 1606 1698
rect 905 1449 910 1487
rect 1007 1445 1012 1463
rect 1601 1440 1606 1522
rect 905 1273 910 1311
rect 1007 1269 1012 1287
rect 1601 1264 1606 1346
rect 905 1097 910 1135
rect 1007 1093 1012 1111
rect 1601 1088 1606 1170
rect 905 921 910 959
rect 1007 917 1012 935
rect 1601 912 1606 994
rect 905 745 910 783
rect 1007 741 1012 759
rect 1601 736 1606 818
rect 905 569 910 607
rect 1007 565 1012 583
rect 1601 560 1606 642
rect 1687 542 1692 1893
rect 1771 1827 1776 1867
rect 1785 1843 1786 1848
rect 1781 1834 1786 1843
rect 1793 1834 1798 1885
rect 1946 1876 1951 1879
rect 2019 1876 2024 1879
rect 2053 1876 2058 1880
rect 2126 1876 2131 1880
rect 2246 1876 2251 1880
rect 2319 1876 2324 1880
rect 1807 1834 1812 1867
rect 1820 1796 1825 1828
rect 2401 1792 2406 1874
rect 2571 1827 2576 1867
rect 2585 1843 2586 1848
rect 2581 1834 2586 1843
rect 2593 1834 2598 1885
rect 2607 1834 2612 1867
rect 2695 1827 2700 1867
rect 2709 1843 2710 1848
rect 2705 1834 2710 1843
rect 2717 1834 2722 1885
rect 2731 1834 2736 1867
rect 2819 1827 2824 1867
rect 2833 1843 2834 1848
rect 2829 1834 2834 1843
rect 2841 1834 2846 1885
rect 2855 1834 2860 1867
rect 2635 1778 2640 1799
rect 2759 1769 2764 1799
rect 1820 1620 1825 1652
rect 2401 1616 2406 1698
rect 2635 1602 2640 1623
rect 2759 1593 2764 1623
rect 1820 1444 1825 1476
rect 2401 1440 2406 1522
rect 2635 1426 2640 1447
rect 2759 1417 2764 1447
rect 1820 1268 1825 1300
rect 2401 1264 2406 1346
rect 2635 1250 2640 1271
rect 2759 1241 2764 1271
rect 1820 1092 1825 1124
rect 2401 1088 2406 1170
rect 2635 1074 2640 1095
rect 2759 1065 2764 1095
rect 1820 916 1825 948
rect 2401 912 2406 994
rect 2635 898 2640 919
rect 2759 889 2764 919
rect 1820 740 1825 772
rect 2401 736 2406 818
rect 2635 722 2640 743
rect 2759 713 2764 743
rect 1820 564 1825 596
rect 2401 560 2406 642
rect 2635 546 2640 567
rect 2759 537 2764 567
<< m234contact >>
rect 164 1893 169 1898
rect 164 1882 169 1887
rect 164 1870 169 1875
rect 47 1810 52 1815
rect 447 1856 452 1861
rect 447 1800 452 1805
rect 437 1793 442 1798
rect 644 1793 649 1798
rect 734 1711 739 1732
rect 447 1680 452 1685
rect 47 1634 52 1639
rect 447 1624 452 1629
rect 437 1617 442 1622
rect 644 1617 649 1622
rect 447 1504 452 1509
rect 47 1458 52 1463
rect 447 1448 452 1453
rect 437 1441 442 1446
rect 644 1441 649 1446
rect 447 1328 452 1333
rect 47 1282 52 1287
rect 447 1272 452 1277
rect 437 1265 442 1270
rect 644 1265 649 1270
rect 447 1152 452 1157
rect 47 1106 52 1111
rect 447 1096 452 1101
rect 437 1089 442 1094
rect 644 1089 649 1094
rect 447 976 452 981
rect 47 930 52 935
rect 447 920 452 925
rect 437 913 442 918
rect 644 913 649 918
rect 447 800 452 805
rect 47 754 52 759
rect 447 744 452 749
rect 437 737 442 742
rect 644 737 649 742
rect 447 624 452 629
rect 47 578 52 583
rect 447 568 452 573
rect 437 561 442 566
rect 644 561 649 566
rect 2521 1893 2526 1898
rect 1338 1850 1343 1855
rect 905 1839 910 1844
rect 1012 1839 1017 1844
rect 1119 1839 1124 1844
rect 1226 1839 1231 1844
rect 905 1796 910 1801
rect 1007 1792 1012 1797
rect 1114 1792 1119 1797
rect 1221 1792 1226 1797
rect 1328 1792 1333 1797
rect 1338 1791 1343 1796
rect 1007 1773 1012 1778
rect 1114 1773 1119 1778
rect 1221 1773 1226 1778
rect 1328 1773 1333 1778
rect 1528 1773 1533 1778
rect 838 1741 843 1762
rect 1551 1741 1556 1760
rect 1609 1711 1614 1732
rect 1338 1674 1343 1679
rect 905 1663 910 1668
rect 1012 1663 1017 1668
rect 1119 1663 1124 1668
rect 1226 1663 1231 1668
rect 905 1620 910 1625
rect 1007 1616 1012 1621
rect 1114 1616 1119 1621
rect 1221 1616 1226 1621
rect 1328 1616 1333 1621
rect 1338 1615 1343 1620
rect 1007 1597 1012 1602
rect 1114 1597 1119 1602
rect 1221 1597 1226 1602
rect 1328 1597 1333 1602
rect 1528 1597 1533 1602
rect 1338 1498 1343 1503
rect 905 1487 910 1492
rect 1012 1487 1017 1492
rect 1119 1487 1124 1492
rect 1226 1487 1231 1492
rect 905 1444 910 1449
rect 1007 1440 1012 1445
rect 1114 1440 1119 1445
rect 1221 1440 1226 1445
rect 1328 1440 1333 1445
rect 1338 1439 1343 1444
rect 1007 1421 1012 1426
rect 1114 1421 1119 1426
rect 1221 1421 1226 1426
rect 1328 1421 1333 1426
rect 1528 1421 1533 1426
rect 1338 1322 1343 1327
rect 905 1311 910 1316
rect 1012 1311 1017 1316
rect 1119 1311 1124 1316
rect 1226 1311 1231 1316
rect 905 1268 910 1273
rect 1007 1264 1012 1269
rect 1114 1264 1119 1269
rect 1221 1264 1226 1269
rect 1328 1264 1333 1269
rect 1338 1263 1343 1268
rect 1007 1245 1012 1250
rect 1114 1245 1119 1250
rect 1221 1245 1226 1250
rect 1328 1245 1333 1250
rect 1528 1245 1533 1250
rect 1338 1146 1343 1151
rect 905 1135 910 1140
rect 1012 1135 1017 1140
rect 1119 1135 1124 1140
rect 1226 1135 1231 1140
rect 905 1092 910 1097
rect 1007 1088 1012 1093
rect 1114 1088 1119 1093
rect 1221 1088 1226 1093
rect 1328 1088 1333 1093
rect 1338 1087 1343 1092
rect 1007 1069 1012 1074
rect 1114 1069 1119 1074
rect 1221 1069 1226 1074
rect 1328 1069 1333 1074
rect 1528 1069 1533 1074
rect 1338 970 1343 975
rect 905 959 910 964
rect 1012 959 1017 964
rect 1119 959 1124 964
rect 1226 959 1231 964
rect 905 916 910 921
rect 1007 912 1012 917
rect 1114 912 1119 917
rect 1221 912 1226 917
rect 1328 912 1333 917
rect 1338 911 1343 916
rect 1007 893 1012 898
rect 1114 893 1119 898
rect 1221 893 1226 898
rect 1328 893 1333 898
rect 1528 893 1533 898
rect 1338 794 1343 799
rect 905 783 910 788
rect 1012 783 1017 788
rect 1119 783 1124 788
rect 1226 783 1231 788
rect 905 740 910 745
rect 1007 736 1012 741
rect 1114 736 1119 741
rect 1221 736 1226 741
rect 1328 736 1333 741
rect 1338 735 1343 740
rect 1007 717 1012 722
rect 1114 717 1119 722
rect 1221 717 1226 722
rect 1328 717 1333 722
rect 1528 717 1533 722
rect 1338 618 1343 623
rect 905 607 910 612
rect 1012 607 1017 612
rect 1119 607 1124 612
rect 1226 607 1231 612
rect 905 564 910 569
rect 1007 560 1012 565
rect 1114 560 1119 565
rect 1221 560 1226 565
rect 1328 560 1333 565
rect 1338 559 1343 564
rect 1007 541 1012 546
rect 1114 541 1119 546
rect 1221 541 1226 546
rect 1328 541 1333 546
rect 1528 541 1533 546
rect 1838 1850 1843 1855
rect 2138 1850 2143 1855
rect 2032 1839 2037 1844
rect 1849 1796 1854 1801
rect 2028 1792 2033 1797
rect 2143 1796 2148 1801
rect 2328 1792 2333 1797
rect 2626 1796 2631 1801
rect 2135 1773 2140 1778
rect 2028 1764 2033 1769
rect 2328 1764 2333 1769
rect 2351 1741 2356 1760
rect 2409 1711 2414 1732
rect 1838 1674 1843 1679
rect 2138 1674 2143 1679
rect 2032 1663 2037 1668
rect 1849 1620 1854 1625
rect 2028 1616 2033 1621
rect 2143 1620 2148 1625
rect 2328 1616 2333 1621
rect 2626 1620 2631 1625
rect 2135 1597 2140 1602
rect 2028 1588 2033 1593
rect 2328 1588 2333 1593
rect 1838 1498 1843 1503
rect 2138 1498 2143 1503
rect 2032 1487 2037 1492
rect 1849 1444 1854 1449
rect 2028 1440 2033 1445
rect 2143 1444 2148 1449
rect 2328 1440 2333 1445
rect 2626 1444 2631 1449
rect 2135 1421 2140 1426
rect 2028 1412 2033 1417
rect 2328 1412 2333 1417
rect 1838 1322 1843 1327
rect 2138 1322 2143 1327
rect 2032 1311 2037 1316
rect 1849 1268 1854 1273
rect 2028 1264 2033 1269
rect 2143 1268 2148 1273
rect 2328 1264 2333 1269
rect 2626 1268 2631 1273
rect 2135 1245 2140 1250
rect 2028 1236 2033 1241
rect 2328 1236 2333 1241
rect 1838 1146 1843 1151
rect 2138 1146 2143 1151
rect 2032 1135 2037 1140
rect 1849 1092 1854 1097
rect 2028 1088 2033 1093
rect 2143 1092 2148 1097
rect 2328 1088 2333 1093
rect 2626 1092 2631 1097
rect 2135 1069 2140 1074
rect 2028 1060 2033 1065
rect 2328 1060 2333 1065
rect 1838 970 1843 975
rect 2138 970 2143 975
rect 2032 959 2037 964
rect 1849 916 1854 921
rect 2028 912 2033 917
rect 2143 916 2148 921
rect 2328 912 2333 917
rect 2626 916 2631 921
rect 2135 893 2140 898
rect 2028 884 2033 889
rect 2328 884 2333 889
rect 1838 794 1843 799
rect 2138 794 2143 799
rect 2032 783 2037 788
rect 1849 740 1854 745
rect 2028 736 2033 741
rect 2143 740 2148 745
rect 2328 736 2333 741
rect 2626 740 2631 745
rect 2135 717 2140 722
rect 2028 708 2033 713
rect 2328 708 2333 713
rect 1838 618 1843 623
rect 2138 618 2143 623
rect 2032 607 2037 612
rect 1849 564 1854 569
rect 2028 560 2033 565
rect 2143 564 2148 569
rect 2328 560 2333 565
rect 2626 564 2631 569
rect 2135 541 2140 546
rect 2028 532 2033 537
rect 2328 532 2333 537
<< m4contact >>
rect 635 1972 640 1977
rect 914 1972 919 1977
rect 635 1882 640 1887
rect 428 1870 433 1875
rect 684 1856 689 1861
rect 165 1793 170 1798
rect 201 1775 206 1780
rect 726 1805 731 1820
rect 38 1770 43 1775
rect 447 1770 452 1775
rect 684 1773 689 1778
rect -42 1741 -37 1762
rect 17 1741 22 1762
rect 68 1741 73 1762
rect 127 1741 132 1762
rect 245 1741 250 1762
rect 391 1741 396 1762
rect 505 1743 510 1770
rect 598 1741 603 1762
rect -30 1711 -25 1732
rect 29 1711 34 1732
rect 56 1711 61 1732
rect 115 1711 120 1732
rect 264 1711 269 1732
rect 379 1711 384 1732
rect 577 1711 582 1732
rect 586 1711 591 1732
rect 684 1680 689 1685
rect 165 1617 170 1622
rect 201 1599 206 1604
rect 726 1629 731 1644
rect 38 1594 43 1599
rect 447 1594 452 1599
rect 684 1597 689 1602
rect 684 1504 689 1509
rect 165 1441 170 1446
rect 201 1423 206 1428
rect 726 1453 731 1468
rect 38 1418 43 1423
rect 447 1418 452 1423
rect 684 1421 689 1426
rect 684 1328 689 1333
rect 165 1265 170 1270
rect 201 1247 206 1252
rect 726 1277 731 1292
rect 38 1242 43 1247
rect 447 1242 452 1247
rect 684 1245 689 1250
rect 684 1152 689 1157
rect 165 1089 170 1094
rect 201 1071 206 1076
rect 726 1101 731 1116
rect 38 1066 43 1071
rect 447 1066 452 1071
rect 684 1069 689 1074
rect 684 976 689 981
rect 165 913 170 918
rect 201 895 206 900
rect 726 925 731 940
rect 38 890 43 895
rect 447 890 452 895
rect 684 893 689 898
rect 684 800 689 805
rect 165 737 170 742
rect 201 719 206 724
rect 726 749 731 764
rect 38 714 43 719
rect 447 714 452 719
rect 684 717 689 722
rect 684 624 689 629
rect 165 561 170 566
rect 201 543 206 548
rect 726 573 731 588
rect 38 538 43 543
rect 447 538 452 543
rect 684 541 689 546
rect 914 1956 919 1961
rect 962 1956 967 1961
rect 896 1893 901 1898
rect 1687 1893 1692 1898
rect 896 1863 901 1868
rect 1007 1815 1012 1820
rect 859 1741 864 1762
rect 952 1741 957 1762
rect 1059 1741 1064 1762
rect 1166 1741 1171 1762
rect 1273 1741 1278 1762
rect 1426 1741 1431 1760
rect 1473 1741 1478 1760
rect 847 1711 852 1732
rect 934 1711 939 1732
rect 1041 1711 1046 1732
rect 1148 1711 1153 1732
rect 1255 1711 1260 1732
rect 1381 1711 1386 1732
rect 1455 1711 1460 1732
rect 1007 1639 1012 1644
rect 1007 1463 1012 1468
rect 1007 1287 1012 1292
rect 1007 1111 1012 1116
rect 1007 935 1012 940
rect 1007 759 1012 764
rect 1007 583 1012 588
rect 1820 1791 1825 1796
rect 2635 1773 2640 1778
rect 2759 1764 2764 1769
rect 1734 1741 1739 1760
rect 1793 1741 1798 1760
rect 1926 1741 1931 1760
rect 1973 1741 1978 1760
rect 2080 1741 2085 1760
rect 2226 1741 2231 1760
rect 2273 1741 2278 1760
rect 2534 1741 2539 1760
rect 2593 1741 2598 1760
rect 2658 1741 2663 1760
rect 2717 1741 2722 1760
rect 2782 1741 2787 1760
rect 2841 1741 2846 1760
rect 1722 1711 1727 1732
rect 1781 1711 1786 1732
rect 1881 1711 1886 1732
rect 1955 1711 1960 1732
rect 2062 1711 2067 1732
rect 2181 1711 2186 1732
rect 2255 1711 2260 1732
rect 2522 1711 2527 1732
rect 2581 1711 2586 1732
rect 2646 1711 2651 1732
rect 2705 1711 2710 1732
rect 2770 1711 2775 1732
rect 2829 1711 2834 1732
rect 1820 1615 1825 1620
rect 2635 1597 2640 1602
rect 2759 1588 2764 1593
rect 1820 1439 1825 1444
rect 2635 1421 2640 1426
rect 2759 1412 2764 1417
rect 1820 1263 1825 1268
rect 2635 1245 2640 1250
rect 2759 1236 2764 1241
rect 1820 1087 1825 1092
rect 2635 1069 2640 1074
rect 2759 1060 2764 1065
rect 1820 911 1825 916
rect 2635 893 2640 898
rect 2759 884 2764 889
rect 1820 735 1825 740
rect 2635 717 2640 722
rect 2759 708 2764 713
rect 1820 559 1825 564
rect 2635 541 2640 546
rect 2759 532 2764 537
<< metal4 >>
rect 640 1972 914 1977
rect 919 1956 962 1961
rect 169 1893 896 1898
rect 1692 1893 2521 1898
rect 169 1882 635 1887
rect 169 1870 428 1875
rect 452 1856 684 1861
rect 1343 1850 1838 1855
rect 1843 1850 2138 1855
rect 1338 1849 1343 1850
rect 1226 1844 1343 1849
rect 2032 1844 2037 1850
rect 910 1839 1012 1844
rect 1017 1839 1119 1844
rect 1124 1839 1226 1844
rect 447 1805 726 1810
rect 731 1815 1007 1820
rect 1849 1801 2631 1806
rect 170 1793 437 1798
rect 905 1793 910 1796
rect 437 1788 910 1793
rect 1012 1792 1114 1797
rect 1119 1792 1221 1797
rect 1226 1792 1328 1797
rect 1343 1791 1820 1796
rect 2028 1787 2333 1792
rect 43 1770 447 1775
rect 689 1773 1007 1778
rect 1012 1773 1114 1778
rect 1119 1773 1221 1778
rect 1226 1773 1328 1778
rect 1333 1773 1528 1778
rect 1533 1773 2135 1778
rect 2140 1773 2635 1778
rect -81 1741 -42 1762
rect -37 1741 17 1762
rect 22 1741 68 1762
rect 73 1741 127 1762
rect 132 1741 245 1762
rect 250 1741 391 1762
rect 396 1743 505 1762
rect 2033 1764 2328 1769
rect 2333 1764 2759 1769
rect 510 1743 598 1762
rect 396 1741 598 1743
rect 603 1741 838 1762
rect 843 1741 859 1762
rect 864 1741 952 1762
rect 957 1741 1059 1762
rect 1064 1741 1166 1762
rect 1171 1741 1273 1762
rect 1278 1760 1324 1762
rect 1278 1741 1426 1760
rect 1431 1741 1473 1760
rect 1478 1741 1551 1760
rect 1556 1741 1734 1760
rect 1739 1741 1793 1760
rect 1798 1741 1926 1760
rect 1931 1741 1973 1760
rect 1978 1741 2080 1760
rect 2085 1741 2226 1760
rect 2231 1741 2273 1760
rect 2278 1741 2351 1760
rect 2356 1741 2534 1760
rect 2539 1741 2593 1760
rect 2598 1741 2658 1760
rect 2663 1741 2717 1760
rect 2722 1741 2782 1760
rect 2787 1741 2841 1760
rect 2846 1741 2885 1760
rect -81 1711 -30 1732
rect -25 1711 29 1732
rect 34 1711 56 1732
rect 61 1711 115 1732
rect 120 1711 264 1732
rect 269 1711 379 1732
rect 384 1711 577 1732
rect 582 1711 586 1732
rect 591 1711 734 1732
rect 739 1711 847 1732
rect 852 1711 934 1732
rect 939 1711 1041 1732
rect 1046 1711 1148 1732
rect 1153 1711 1255 1732
rect 1260 1711 1381 1732
rect 1386 1711 1455 1732
rect 1460 1711 1609 1732
rect 1614 1711 1722 1732
rect 1727 1711 1781 1732
rect 1786 1711 1881 1732
rect 1886 1711 1955 1732
rect 1960 1711 2062 1732
rect 2067 1711 2181 1732
rect 2186 1711 2255 1732
rect 2260 1711 2409 1732
rect 2414 1711 2522 1732
rect 2527 1711 2581 1732
rect 2586 1711 2646 1732
rect 2651 1711 2705 1732
rect 2710 1711 2770 1732
rect 2775 1711 2829 1732
rect 2834 1711 2885 1732
rect 452 1680 684 1685
rect 1343 1674 1838 1679
rect 1843 1674 2138 1679
rect 1338 1673 1343 1674
rect 1226 1668 1343 1673
rect 2032 1668 2037 1674
rect 910 1663 1012 1668
rect 1017 1663 1119 1668
rect 1124 1663 1226 1668
rect 447 1629 726 1634
rect 731 1639 1007 1644
rect 1849 1625 2631 1630
rect 170 1617 437 1622
rect 905 1617 910 1620
rect 437 1612 910 1617
rect 1012 1616 1114 1621
rect 1119 1616 1221 1621
rect 1226 1616 1328 1621
rect 1343 1615 1820 1620
rect 2028 1611 2333 1616
rect 43 1594 447 1599
rect 689 1597 1007 1602
rect 1012 1597 1114 1602
rect 1119 1597 1221 1602
rect 1226 1597 1328 1602
rect 1333 1597 1528 1602
rect 1533 1597 2135 1602
rect 2140 1597 2635 1602
rect 2033 1588 2328 1593
rect 2333 1588 2759 1593
rect 452 1504 684 1509
rect 1343 1498 1838 1503
rect 1843 1498 2138 1503
rect 1338 1497 1343 1498
rect 1226 1492 1343 1497
rect 2032 1492 2037 1498
rect 910 1487 1012 1492
rect 1017 1487 1119 1492
rect 1124 1487 1226 1492
rect 447 1453 726 1458
rect 731 1463 1007 1468
rect 1849 1449 2631 1454
rect 170 1441 437 1446
rect 905 1441 910 1444
rect 437 1436 910 1441
rect 1012 1440 1114 1445
rect 1119 1440 1221 1445
rect 1226 1440 1328 1445
rect 1343 1439 1820 1444
rect 2028 1435 2333 1440
rect 43 1418 447 1423
rect 689 1421 1007 1426
rect 1012 1421 1114 1426
rect 1119 1421 1221 1426
rect 1226 1421 1328 1426
rect 1333 1421 1528 1426
rect 1533 1421 2135 1426
rect 2140 1421 2635 1426
rect 2033 1412 2328 1417
rect 2333 1412 2759 1417
rect 452 1328 684 1333
rect 1343 1322 1838 1327
rect 1843 1322 2138 1327
rect 1338 1321 1343 1322
rect 1226 1316 1343 1321
rect 2032 1316 2037 1322
rect 910 1311 1012 1316
rect 1017 1311 1119 1316
rect 1124 1311 1226 1316
rect 447 1277 726 1282
rect 731 1287 1007 1292
rect 1849 1273 2631 1278
rect 170 1265 437 1270
rect 905 1265 910 1268
rect 437 1260 910 1265
rect 1012 1264 1114 1269
rect 1119 1264 1221 1269
rect 1226 1264 1328 1269
rect 1343 1263 1820 1268
rect 2028 1259 2333 1264
rect 43 1242 447 1247
rect 689 1245 1007 1250
rect 1012 1245 1114 1250
rect 1119 1245 1221 1250
rect 1226 1245 1328 1250
rect 1333 1245 1528 1250
rect 1533 1245 2135 1250
rect 2140 1245 2635 1250
rect 2033 1236 2328 1241
rect 2333 1236 2759 1241
rect 452 1152 684 1157
rect 1343 1146 1838 1151
rect 1843 1146 2138 1151
rect 1338 1145 1343 1146
rect 1226 1140 1343 1145
rect 2032 1140 2037 1146
rect 910 1135 1012 1140
rect 1017 1135 1119 1140
rect 1124 1135 1226 1140
rect 447 1101 726 1106
rect 731 1111 1007 1116
rect 1849 1097 2631 1102
rect 170 1089 437 1094
rect 905 1089 910 1092
rect 437 1084 910 1089
rect 1012 1088 1114 1093
rect 1119 1088 1221 1093
rect 1226 1088 1328 1093
rect 1343 1087 1820 1092
rect 2028 1083 2333 1088
rect 43 1066 447 1071
rect 689 1069 1007 1074
rect 1012 1069 1114 1074
rect 1119 1069 1221 1074
rect 1226 1069 1328 1074
rect 1333 1069 1528 1074
rect 1533 1069 2135 1074
rect 2140 1069 2635 1074
rect 2033 1060 2328 1065
rect 2333 1060 2759 1065
rect 452 976 684 981
rect 1343 970 1838 975
rect 1843 970 2138 975
rect 1338 969 1343 970
rect 1226 964 1343 969
rect 2032 964 2037 970
rect 910 959 1012 964
rect 1017 959 1119 964
rect 1124 959 1226 964
rect 447 925 726 930
rect 731 935 1007 940
rect 1849 921 2631 926
rect 170 913 437 918
rect 905 913 910 916
rect 437 908 910 913
rect 1012 912 1114 917
rect 1119 912 1221 917
rect 1226 912 1328 917
rect 1343 911 1820 916
rect 2028 907 2333 912
rect 43 890 447 895
rect 689 893 1007 898
rect 1012 893 1114 898
rect 1119 893 1221 898
rect 1226 893 1328 898
rect 1333 893 1528 898
rect 1533 893 2135 898
rect 2140 893 2635 898
rect 2033 884 2328 889
rect 2333 884 2759 889
rect 452 800 684 805
rect 1343 794 1838 799
rect 1843 794 2138 799
rect 1338 793 1343 794
rect 1226 788 1343 793
rect 2032 788 2037 794
rect 910 783 1012 788
rect 1017 783 1119 788
rect 1124 783 1226 788
rect 447 749 726 754
rect 731 759 1007 764
rect 1849 745 2631 750
rect 170 737 437 742
rect 905 737 910 740
rect 437 732 910 737
rect 1012 736 1114 741
rect 1119 736 1221 741
rect 1226 736 1328 741
rect 1343 735 1820 740
rect 2028 731 2333 736
rect 43 714 447 719
rect 689 717 1007 722
rect 1012 717 1114 722
rect 1119 717 1221 722
rect 1226 717 1328 722
rect 1333 717 1528 722
rect 1533 717 2135 722
rect 2140 717 2635 722
rect 2033 708 2328 713
rect 2333 708 2759 713
rect 452 624 684 629
rect 1343 618 1838 623
rect 1843 618 2138 623
rect 1338 617 1343 618
rect 1226 612 1343 617
rect 2032 612 2037 618
rect 910 607 1012 612
rect 1017 607 1119 612
rect 1124 607 1226 612
rect 447 573 726 578
rect 731 583 1007 588
rect 1849 569 2631 574
rect 170 561 437 566
rect 905 561 910 564
rect 437 556 910 561
rect 1012 560 1114 565
rect 1119 560 1221 565
rect 1226 560 1328 565
rect 1343 559 1820 564
rect 2028 555 2333 560
rect 43 538 447 543
rect 689 541 1007 546
rect 1012 541 1114 546
rect 1119 541 1221 546
rect 1226 541 1328 546
rect 1333 541 1528 546
rect 1533 541 2135 546
rect 2140 541 2635 546
rect 2033 532 2328 537
rect 2333 532 2759 537
use staticizer  staticizer_1
timestamp 1765745113
transform -1 0 39 0 1 1753
box 61 -1215 120 78
use latch  latch_4
timestamp 1765416915
transform -1 0 -355 0 1 463
box -392 82 -333 1369
use latch  latch_0
timestamp 1765416915
transform 1 0 445 0 1 463
box -392 82 -333 1369
use 4nor2  4nor2_0
timestamp 1761285742
transform 0 1 81 -1 0 1980
box 68 -24 135 80
use inv2  inv2_0
timestamp 1765338958
transform -1 0 -22 0 1 1852
box -10 -13 20 40
use staticizer  staticizer_0
timestamp 1765745113
transform 1 0 51 0 1 1753
box 61 -1215 120 78
use shift  shift_0
timestamp 1765416915
transform 1 0 330 0 1 2153
box -138 -1615 46 -268
use latch  latch_3
timestamp 1765416915
transform 1 0 768 0 1 456
box -392 82 -333 1369
use fblock  fblock_0
timestamp 1765416915
transform 1 0 535 0 1 2993
box -80 -2455 50 -1047
use latch  latch_1
timestamp 1765416915
transform 1 0 975 0 1 456
box -392 82 -333 1369
use addsub  addsub_0
timestamp 1765338694
transform 1 0 675 0 1 712
box -14 -174 166 1225
use staticizer_one  staticizer_one_0
timestamp 1765328088
transform 1 0 867 0 1 1967
box 54 -61 113 -1
use latch  latch_2
timestamp 1765416915
transform 1 0 1236 0 1 459
box -392 82 -333 1369
use reg  reg_0
timestamp 1765316199
transform 1 0 928 0 1 936
box -14 -398 76 940
use reg  reg_1
timestamp 1765316199
transform 1 0 1035 0 1 936
box -14 -398 76 940
use 2nor  2nor_0
timestamp 1762488699
transform -1 0 1042 0 1 1940
box 68 28 115 81
use latch_one  latch_one_1
timestamp 1765002978
transform 1 0 873 0 1 2033
box -11 -67 48 -12
use reg_one  reg_one_0
timestamp 1761015633
transform 1 0 991 0 1 1924
box -11 -25 74 81
use latch_one  latch_one_0
timestamp 1765002978
transform 1 0 873 0 1 1978
box -11 -67 48 -12
use reg  reg_2
timestamp 1765316199
transform 1 0 1142 0 1 936
box -14 -398 76 940
use mux_8bit  mux_8bit_0
timestamp 1765349323
transform 1 0 1342 0 1 1766
box 1 -1228 92 116
use reg  reg_3
timestamp 1765316199
transform 1 0 1249 0 1 936
box -14 -398 76 940
use inv2  inv2_6
timestamp 1765338958
transform 0 -1 1417 -1 0 1926
box -10 -13 20 40
use inv2  inv2_3
timestamp 1765338958
transform 0 -1 1417 -1 0 1896
box -10 -13 20 40
use inv2  inv2_8
timestamp 1765338958
transform 0 -1 1417 -1 0 1986
box -10 -13 20 40
use inv2  inv2_7
timestamp 1765338958
transform 0 -1 1417 -1 0 1956
box -10 -13 20 40
use addsub  addsub_1
timestamp 1765338694
transform 1 0 1550 0 1 712
box -14 -174 166 1225
use reg  reg_4
timestamp 1765316199
transform 1 0 1449 0 1 936
box -14 -398 76 940
use latch  latch_5
timestamp 1765416915
transform 1 0 2111 0 1 459
box -392 82 -333 1369
use inv2  inv2_4
timestamp 1765338958
transform 1 0 1776 0 -1 1880
box -10 -13 20 40
use staticizer  staticizer_2
timestamp 1765745113
transform 1 0 1717 0 1 1756
box 61 -1215 120 78
use reg  reg_5
timestamp 1765316199
transform 1 0 1949 0 1 936
box -14 -398 76 940
use mux_8bit  mux_8bit_1
timestamp 1765349323
transform 1 0 1842 0 1 1766
box 1 -1228 92 116
use inv2  inv2_12
timestamp 1765338958
transform 0 -1 1917 -1 0 1926
box -10 -13 20 40
use inv2  inv2_11
timestamp 1765338958
transform 0 -1 1917 -1 0 1896
box -10 -13 20 40
use inv2  inv2_10
timestamp 1765338958
transform 0 -1 1917 -1 0 1956
box -10 -13 20 40
use inv2  inv2_9
timestamp 1765338958
transform 0 -1 1917 -1 0 1986
box -10 -13 20 40
use reg  reg_6
timestamp 1765316199
transform 1 0 2056 0 1 936
box -14 -398 76 940
use mux_8bit  mux_8bit_2
timestamp 1765349323
transform 1 0 2142 0 1 1766
box 1 -1228 92 116
use reg  reg_7
timestamp 1765316199
transform 1 0 2249 0 1 936
box -14 -398 76 940
use inv2  inv2_16
timestamp 1765338958
transform 0 -1 2217 -1 0 1926
box -10 -13 20 40
use inv2  inv2_15
timestamp 1765338958
transform 0 -1 2217 -1 0 1896
box -10 -13 20 40
use inv2  inv2_14
timestamp 1765338958
transform 0 -1 2217 -1 0 1986
box -10 -13 20 40
use inv2  inv2_13
timestamp 1765338958
transform 0 -1 2217 -1 0 1956
box -10 -13 20 40
use addsub  addsub_2
timestamp 1765338694
transform 1 0 2350 0 1 712
box -14 -174 166 1225
use staticizer  staticizer_3
timestamp 1765745113
transform 1 0 2517 0 1 1756
box 61 -1215 120 78
use latch  latch_7
timestamp 1765416915
transform 1 0 3035 0 1 459
box -392 82 -333 1369
use latch  latch_6
timestamp 1765416915
transform 1 0 2911 0 1 459
box -392 82 -333 1369
use inv2  inv2_5
timestamp 1765338958
transform 1 0 2576 0 -1 1880
box -10 -13 20 40
use inv2  inv2_1
timestamp 1765338958
transform 1 0 2700 0 -1 1880
box -10 -13 20 40
use staticizer  staticizer_5
timestamp 1765745113
transform 1 0 2765 0 1 1756
box 61 -1215 120 78
use staticizer  staticizer_4
timestamp 1765745113
transform 1 0 2641 0 1 1756
box 61 -1215 120 78
use latch  latch_8
timestamp 1765416915
transform 1 0 3159 0 1 459
box -392 82 -333 1369
use inv2  inv2_2
timestamp 1765338958
transform 1 0 2824 0 -1 1880
box -10 -13 20 40
<< labels >>
rlabel m234contact 47 1810 52 1815 1 data_in0
rlabel m234contact 47 1634 52 1639 1 data_in1
rlabel m234contact 47 1458 52 1463 1 data_in2
rlabel m234contact 47 1282 52 1287 1 data_in3
rlabel m234contact 47 1106 52 1111 1 data_in4
rlabel m234contact 47 930 52 935 1 data_in5
rlabel m234contact 47 754 52 759 1 data_in6
rlabel m234contact 47 578 52 583 1 data_in7
rlabel metal1 -80 1825 -75 1830 3 data_out0
rlabel metal1 -80 1649 -75 1654 3 data_out1
rlabel metal1 -80 1473 -75 1478 3 data_out2
rlabel metal1 -80 1297 -75 1302 3 data_out3
rlabel metal1 -80 1121 -75 1126 3 data_out4
rlabel metal1 -80 945 -75 950 3 data_out5
rlabel metal1 -80 769 -75 774 3 data_out6
rlabel metal1 -80 593 -75 598 3 data_out7
rlabel metal3 284 1885 289 1887 1 os_u
rlabel metal3 346 1885 351 1887 1 os_s
rlabel metal3 428 1824 433 1828 1 ros
rlabel metal3 456 1922 461 1948 1 fb_g3
rlabel metal3 488 1922 493 1948 1 fb_g2
rlabel metal3 522 1922 527 1948 1 fb_g1
rlabel metal3 555 1922 560 1948 1 fb_g0
rlabel metal3 635 1824 640 1828 1 rfb
rlabel metal1 812 538 817 543 1 as_cout
rlabel metal1 661 1829 666 1834 1 as_sub
rlabel metal1 842 1898 847 1901 1 as_cin
rlabel metal2 914 1876 919 1880 1 A_r0
rlabel metal3 925 1876 930 1880 1 A_r1
rlabel metal3 998 1876 1003 1880 1 A_w
rlabel metal2 1021 1876 1026 1880 1 DB_r0
rlabel metal3 1032 1876 1037 1880 1 DB_r1
rlabel metal3 1105 1876 1110 1880 1 DB_w
rlabel metal3 1139 1876 1144 1880 1 X_r1
rlabel metal2 1128 1876 1133 1880 1 X_r0
rlabel metal3 1212 1876 1217 1880 1 X_w
rlabel metal2 1235 1876 1240 1880 1 Y_r0
rlabel metal3 1246 1876 1251 1880 1 Y_r1
rlabel metal3 1319 1876 1324 1880 1 Y_w
rlabel metal3 1446 1876 1451 1879 1 PCL_r1
rlabel metal3 1519 1876 1524 1879 1 PCL_w
rlabel metal2 1435 1876 1440 1879 1 PCL_r0
rlabel metal3 1771 1835 1776 1838 1 rPCplus1L
rlabel metal3 2571 1834 2576 1838 1 rPCplus1H
rlabel metal3 2695 1836 2700 1839 1 rd_addrL
rlabel metal3 2819 1834 2824 1837 1 rd_addrH
rlabel metal2 1935 1876 1940 1879 1 PCH_r0
rlabel metal3 2019 1876 2024 1879 1 PCH_w
rlabel metal3 1946 1876 1951 1879 1 PCH_r1
rlabel metal2 2042 1876 2047 1880 1 ABL_r0
rlabel metal3 2053 1876 2058 1880 1 ABL_r1
rlabel metal3 2126 1876 2131 1880 1 ABL_w
rlabel metal2 2235 1876 2240 1880 1 ABH_r0
rlabel metal3 2246 1876 2251 1880 1 ABH_r1
rlabel metal3 2319 1876 2324 1880 1 ABH_w
rlabel m4contact 38 538 43 543 1 rx7
rlabel m4contact 38 714 43 719 1 rx6
rlabel m4contact 38 890 43 895 1 rx5
rlabel m4contact 38 1066 43 1071 1 rx4
rlabel m4contact 38 1242 43 1247 1 rx3
rlabel m4contact 38 1418 43 1423 1 rx2
rlabel m4contact 38 1770 43 1775 1 rx0
rlabel m4contact 38 1594 43 1599 1 rx1
rlabel m123contact 160 1825 165 1830 1 wz0
rlabel m123contact 160 1649 165 1654 1 wz1
rlabel m123contact 160 1473 165 1478 1 wz2
rlabel m123contact 160 1297 165 1302 1 wz3
rlabel m123contact 160 945 165 950 1 wz5
rlabel m123contact 160 769 165 774 1 wz6
rlabel m123contact 160 593 165 598 1 wz7
rlabel m123contact 160 1121 165 1126 1 wz4
rlabel m234contact 447 1856 452 1861 1 ry0
rlabel m234contact 447 1680 452 1685 1 ry1
rlabel m234contact 447 1504 452 1509 1 ry2
rlabel m234contact 447 1328 452 1333 1 ry3
rlabel m234contact 447 1152 452 1157 1 ry4
rlabel m234contact 447 976 452 981 1 ry5
rlabel m234contact 447 800 452 805 1 ry6
rlabel m234contact 447 624 452 629 1 ry7
rlabel metal4 -81 1741 -75 1762 3 GND!
rlabel metal4 -81 1711 -75 1732 3 Vdd!
rlabel m234contact 1338 1791 1343 1796 1 wz_addrL0
rlabel m234contact 1338 1615 1343 1620 1 wz_addrL1
rlabel m234contact 1338 1439 1343 1444 1 wz_addrL2
rlabel m234contact 1338 1263 1343 1268 1 wz_addrL3
rlabel m234contact 1338 1087 1343 1092 1 wz_addrL4
rlabel m234contact 1338 911 1343 916 1 wz_addrL5
rlabel m234contact 1338 735 1343 740 1 wz_addrL6
rlabel m234contact 1338 559 1343 564 1 wz_addrL7
rlabel m234contact 2028 1764 2033 1769 1 ry_addrH0
rlabel m234contact 2028 1588 2033 1593 1 ry_addrH1
rlabel m234contact 2028 1412 2033 1417 1 ry_addrH2
rlabel m234contact 2028 1236 2033 1241 1 ry_addrH3
rlabel m234contact 2028 1060 2033 1065 1 ry_addrH4
rlabel m234contact 2028 884 2033 889 1 ry_addrH5
rlabel m234contact 2028 708 2033 713 1 ry_addrH6
rlabel m234contact 2028 532 2033 537 1 ry_addrH7
rlabel metal1 2823 1799 2828 1804 1 addr_out8
rlabel metal1 2823 1623 2828 1628 1 addr_out9
rlabel metal1 2823 1447 2828 1452 1 addr_out10
rlabel metal1 2823 1271 2828 1276 1 addr_out11
rlabel metal1 2823 1095 2828 1100 1 addr_out12
rlabel metal1 2823 919 2828 924 1 addr_out13
rlabel metal1 2823 743 2828 748 1 addr_out14
rlabel metal1 2823 567 2828 572 1 addr_out15
rlabel metal1 2699 1800 2704 1804 1 addr_out0
rlabel metal1 2699 1624 2704 1628 1 addr_out1
rlabel metal1 2699 1448 2704 1452 1 addr_out2
rlabel metal1 2699 1272 2704 1276 1 addr_out3
rlabel metal1 2699 1096 2704 1100 1 addr_out4
rlabel metal1 2699 920 2704 924 1 addr_out5
rlabel metal1 2699 744 2704 748 1 addr_out6
rlabel metal1 2699 568 2704 572 1 addr_out7
rlabel metal4 1849 1801 1854 1806 1 wz_addrH0
rlabel metal4 1849 1625 1854 1630 1 wz_addrH1
rlabel metal4 1849 1449 1854 1454 1 wz_addrH2
rlabel metal4 1849 1273 1854 1278 1 wz_addrH3
rlabel metal4 1849 1097 1854 1102 1 wz_addrH4
rlabel metal4 1849 921 1854 926 1 wz_addrH5
rlabel metal4 1849 745 1854 750 1 wz_addrH6
rlabel metal4 1849 569 1854 574 1 wz_addrH7
rlabel m234contact 2028 1792 2033 1797 1 rx_addrH0
rlabel m234contact 2028 1616 2033 1621 1 rx_addrH1
rlabel m234contact 2028 1440 2033 1445 1 rx_addrH2
rlabel m234contact 2028 1264 2033 1269 1 rx_addrH3
rlabel m234contact 2028 1088 2033 1093 1 rx_addrH4
rlabel m234contact 2028 912 2033 917 1 rx_addrH5
rlabel m234contact 2028 736 2033 741 1 rx_addrH6
rlabel m234contact 2028 560 2033 565 1 rx_addrH7
rlabel m2contact 1527 1611 1532 1614 1 rx_PCL1
rlabel m2contact 1527 1435 1532 1438 1 rx_PCL2
rlabel m2contact 1527 1259 1532 1262 1 rx_PCL3
rlabel m2contact 1527 1083 1532 1086 1 rx_PCL4
rlabel m2contact 1527 907 1532 910 1 rx_PCL5
rlabel m2contact 1527 731 1532 734 1 rx_PCL6
rlabel m2contact 1527 555 1532 558 1 rx_PCL7
rlabel m2contact 1527 1787 1532 1790 1 rx_PCL0
rlabel metal3 105 1831 110 1835 1 ld_datain
rlabel metal3 -20 1831 -15 1835 1 rd_dataout
rlabel metal1 1438 1820 1443 1825 1 PCL_w_muxout0
rlabel metal1 1438 1468 1443 1473 1 PCL_w_muxout2
rlabel metal1 1438 1292 1443 1297 1 PCL_w_muxout3
rlabel metal1 1438 1116 1443 1121 1 PCL_w_muxout4
rlabel metal1 1438 940 1443 945 1 PCL_w_muxout5
rlabel metal1 1438 764 1443 769 1 PCL_w_muxout6
rlabel metal1 1438 588 1443 593 1 PCL_w_muxout7
rlabel metal1 1438 1644 1443 1649 1 PCL_w_muxout1
rlabel metal2 1492 1844 1496 1849 1 PCL0
rlabel metal2 1492 1668 1496 1673 1 PCL1
rlabel metal2 1492 1492 1496 1497 1 PCL2
rlabel metal2 1492 1316 1496 1321 1 PCL3
rlabel metal2 1492 1140 1496 1145 1 PCL4
rlabel metal2 1492 964 1496 969 1 PCL5
rlabel metal2 1492 788 1496 793 1 PCL6
rlabel metal2 1492 612 1496 617 1 PCL7
rlabel metal1 1404 1990 1409 1996 5 PCL_w_sel
rlabel metal1 1904 1990 1909 1996 5 PCH_w_sel
rlabel metal1 2204 1991 2209 1996 5 ABH_w_sel
rlabel metal2 1704 1625 1708 1630 1 PCLplus1_1
rlabel metal2 1704 1449 1708 1454 1 PCLplus1_2
rlabel metal2 1704 1273 1708 1278 1 PCLplus1_3
rlabel metal2 1704 1097 1708 1102 1 PCLplus1_4
rlabel metal2 1704 921 1708 926 1 PCLplus1_5
rlabel metal2 1704 745 1708 750 1 PCLplus1_6
rlabel metal2 1704 569 1708 574 1 PCLplus1_7
rlabel metal2 1704 1801 1708 1806 1 PCLplus1_0
rlabel polysilicon 1619 1865 1621 1867 1 addsub1_a0
rlabel metal3 896 1827 901 1833 1 ras
rlabel metal3 1059 2000 1064 2005 5 Cflag_w
rlabel metal2 1058 1902 1063 1907 1 Cflag
<< end >>
