magic
tech scmos
timestamp 1765748214
<< nwell >>
rect -9 -47 40 -18
<< pwell >>
rect -9 -71 40 -48
<< ntransistor >>
rect 4 -59 6 -54
rect 15 -59 17 -54
rect 26 -59 28 -54
<< ptransistor >>
rect 4 -40 6 -30
rect 15 -40 17 -30
rect 26 -40 28 -30
<< ndiffusion >>
rect 2 -59 4 -54
rect 6 -59 15 -54
rect 17 -59 26 -54
rect 28 -59 29 -54
<< pdiffusion >>
rect 2 -40 4 -30
rect 6 -40 8 -30
rect 13 -40 15 -30
rect 17 -40 19 -30
rect 24 -40 26 -30
rect 28 -40 29 -30
<< ndcontact >>
rect -3 -59 2 -54
rect 29 -59 34 -54
<< pdcontact >>
rect -3 -40 2 -30
rect 8 -40 13 -30
rect 19 -40 24 -30
rect 29 -40 34 -30
<< psubstratepcontact >>
rect 19 -68 24 -63
<< nsubstratencontact >>
rect 19 -26 24 -21
<< polysilicon >>
rect 4 -30 6 -27
rect 15 -30 17 -27
rect 26 -30 28 -27
rect 4 -54 6 -40
rect 15 -54 17 -40
rect 26 -54 28 -40
rect 4 -62 6 -59
rect 15 -62 17 -59
rect 26 -62 28 -59
<< metal1 >>
rect -3 -26 19 -21
rect 24 -26 40 -21
rect -3 -30 2 -26
rect 19 -30 24 -26
rect 8 -45 13 -40
rect 29 -45 34 -40
rect 8 -50 40 -45
rect 29 -54 34 -50
rect -3 -63 2 -59
rect -3 -68 19 -63
rect 24 -68 40 -63
<< labels >>
rlabel polysilicon 4 -29 6 -27 1 a
rlabel metal1 35 -68 40 -63 7 GND!
rlabel metal1 35 -26 40 -21 7 Vdd!
rlabel metal1 35 -50 40 -45 7 out
rlabel polysilicon 26 -29 28 -27 1 c
rlabel polysilicon 15 -29 17 -27 1 b
<< end >>
