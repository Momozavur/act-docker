magic
tech scmos
timestamp 1759371655
<< nwell >>
rect 55 -19 122 17
<< pwell >>
rect 55 -54 122 -19
<< ntransistor >>
rect 68 -31 70 -26
rect 87 -31 89 -26
rect 68 -41 70 -36
rect 77 -41 79 -36
rect 98 -41 100 -36
rect 107 -41 109 -36
<< ptransistor >>
rect 68 -1 70 4
rect 77 -1 79 4
rect 98 -1 100 4
rect 107 -1 109 4
rect 68 -11 70 -6
rect 87 -11 89 -6
<< ndiffusion >>
rect 66 -31 68 -26
rect 70 -31 71 -26
rect 86 -31 87 -26
rect 89 -31 91 -26
rect 66 -41 68 -36
rect 70 -41 77 -36
rect 79 -41 91 -36
rect 96 -41 98 -36
rect 100 -41 107 -36
rect 109 -41 111 -36
<< pdiffusion >>
rect 66 -1 68 4
rect 70 -1 71 4
rect 76 -1 77 4
rect 79 -1 81 4
rect 96 -1 98 4
rect 100 -1 107 4
rect 109 -1 111 4
rect 66 -11 68 -6
rect 70 -11 71 -6
rect 86 -11 87 -6
rect 89 -11 91 -6
<< ndcontact >>
rect 71 -31 76 -26
rect 81 -31 86 -26
rect 91 -31 96 -26
rect 61 -41 66 -36
rect 91 -41 96 -36
rect 111 -41 116 -36
<< pdcontact >>
rect 71 -1 76 4
rect 91 -1 96 4
rect 111 -1 116 4
rect 71 -11 76 -6
rect 81 -11 86 -6
rect 91 -11 96 -6
rect 101 -6 106 -1
<< psubstratepcontact >>
rect 91 -51 96 -46
<< nsubstratencontact >>
rect 71 9 76 14
<< polysilicon >>
rect 68 4 70 7
rect 77 4 79 7
rect 98 4 100 7
rect 107 4 109 7
rect 68 -6 70 -1
rect 68 -26 70 -11
rect 68 -36 70 -31
rect 77 -33 79 -1
rect 87 -6 89 -3
rect 87 -26 89 -11
rect 87 -33 89 -31
rect 77 -35 89 -33
rect 77 -36 79 -35
rect 98 -36 100 -1
rect 107 -36 109 -1
rect 68 -44 70 -41
rect 77 -44 79 -41
rect 98 -44 100 -41
rect 107 -44 109 -41
<< polycontact >>
rect 93 -21 98 -16
<< metal1 >>
rect 71 4 76 9
rect 81 4 116 9
rect 71 -6 76 -1
rect 76 -11 81 -6
rect 91 -16 96 -11
rect 91 -21 93 -16
rect 91 -26 96 -21
rect 61 -46 66 -41
rect 76 -46 81 -26
rect 101 -36 106 -6
rect 96 -41 106 -36
rect 111 -46 116 -41
rect 61 -51 91 -46
rect 96 -51 116 -46
<< pm12contact >>
rect 109 -21 114 -16
<< pdm12contact >>
rect 61 -1 66 4
rect 81 -1 86 4
rect 61 -11 66 -6
<< ndm12contact >>
rect 61 -31 66 -26
<< metal2 >>
rect 66 -1 81 4
rect 61 -16 66 -11
rect 61 -21 109 -16
rect 61 -26 66 -21
<< labels >>
rlabel polysilicon 68 -15 70 -13 1 a
rlabel polysilicon 77 -15 79 -13 1 b
rlabel metal1 101 -31 106 -26 1 out
rlabel nsubstratencontact 71 9 76 14 5 Vdd!
rlabel psubstratepcontact 91 -51 96 -46 1 GND!
<< end >>
