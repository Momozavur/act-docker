magic
tech scmos
timestamp 1765766491
<< metal5 >>
rect 10 36 30 40
rect 10 28 14 36
rect 26 28 30 36
rect 10 24 30 28
rect 34 36 56 40
rect 34 28 38 36
rect 52 28 56 36
rect 34 24 56 28
rect 60 36 82 40
rect 60 28 64 36
rect 78 28 82 36
rect 60 24 82 28
rect 10 10 14 24
rect 34 20 46 24
rect 34 10 38 20
rect 42 16 50 20
rect 46 12 54 16
rect 50 10 54 12
rect 60 10 64 24
rect 78 10 82 24
rect 86 36 100 40
rect 108 36 112 40
rect 126 36 130 40
rect 86 14 90 36
rect 96 32 104 36
rect 108 32 116 36
rect 122 32 130 36
rect 100 18 104 32
rect 112 28 126 32
rect 96 14 104 18
rect 86 10 100 14
rect 117 10 121 28
rect 134 14 138 40
rect 152 14 156 40
rect 134 10 156 14
rect 160 36 164 40
rect 160 32 168 36
rect 160 28 172 32
rect 160 10 164 28
rect 168 24 174 28
rect 178 24 182 40
rect 170 20 182 24
rect 176 16 182 20
rect 178 10 182 16
<< end >>
