magic
tech scmos
timestamp 1763591700
<< nwell >>
rect 85 17 227 69
<< pwell >>
rect 85 -15 227 17
<< ntransistor >>
rect 97 -9 99 11
rect 115 -9 117 11
rect 125 -9 127 11
rect 134 -9 136 11
rect 152 -9 154 11
rect 161 -9 163 11
rect 170 -9 172 11
rect 195 -9 197 11
rect 213 -9 215 11
<< ptransistor >>
rect 97 23 99 63
rect 115 23 117 63
rect 125 23 127 63
rect 134 23 136 63
rect 152 23 154 63
rect 161 23 163 63
rect 170 23 172 63
rect 195 23 197 63
rect 213 23 215 63
<< ndiffusion >>
rect 96 -9 97 11
rect 99 -9 100 11
rect 114 -9 115 11
rect 117 -9 118 11
rect 124 -9 125 11
rect 127 -9 128 11
rect 133 -9 134 11
rect 136 -9 137 11
rect 151 -9 152 11
rect 154 -9 161 11
rect 163 -9 164 11
rect 169 -9 170 11
rect 172 -9 173 11
rect 194 -9 195 11
rect 197 -9 198 11
rect 212 -9 213 11
rect 215 -9 216 11
<< pdiffusion >>
rect 96 23 97 63
rect 99 23 100 63
rect 114 23 115 63
rect 117 23 118 63
rect 124 23 125 63
rect 127 23 134 63
rect 136 23 137 63
rect 151 23 152 63
rect 154 23 155 63
rect 160 23 161 63
rect 163 23 164 63
rect 169 23 170 63
rect 172 23 173 63
rect 194 23 195 63
rect 197 23 198 63
rect 212 23 213 63
rect 215 23 216 63
<< ndcontact >>
rect 100 -9 105 11
rect 109 -9 114 11
rect 128 -9 133 11
rect 146 -9 151 11
rect 173 -9 178 11
rect 198 -9 203 11
rect 216 -9 221 11
<< pdcontact >>
rect 100 23 105 63
rect 109 23 114 63
rect 137 23 142 63
rect 155 23 160 63
rect 173 23 178 63
rect 198 23 203 63
rect 216 23 221 63
<< psubstratepdiff >>
rect 187 -9 189 11
<< nsubstratendiff >>
rect 187 23 189 63
<< polysilicon >>
rect 97 63 99 72
rect 115 65 127 67
rect 115 63 117 65
rect 125 63 127 65
rect 134 66 154 68
rect 134 63 136 66
rect 152 63 154 66
rect 161 63 163 72
rect 170 63 172 66
rect 195 63 197 66
rect 213 63 215 66
rect 97 11 99 23
rect 115 18 117 23
rect 108 15 117 18
rect 115 11 117 15
rect 125 11 127 23
rect 134 11 136 23
rect 152 11 154 23
rect 161 11 163 23
rect 170 20 172 23
rect 170 11 172 14
rect 195 11 197 23
rect 213 11 215 23
rect 97 -12 99 -9
rect 115 -12 117 -9
rect 125 -12 127 -9
rect 134 -11 136 -9
rect 152 -11 154 -9
rect 134 -13 154 -11
rect 161 -12 163 -9
rect 170 -12 172 -9
rect 195 -12 197 -9
rect 213 -12 215 -9
rect 143 -18 145 -13
<< polycontact >>
rect 94 72 99 77
rect 158 72 163 77
rect 167 66 172 71
rect 192 66 197 71
rect 103 14 108 19
rect 208 15 213 20
rect 94 -17 99 -12
rect 167 -17 172 -12
rect 142 -23 147 -18
<< metal1 >>
rect 91 72 94 77
rect 133 72 158 75
rect 133 69 136 72
rect 189 71 197 77
rect 111 66 136 69
rect 139 66 167 69
rect 189 69 192 71
rect 175 66 192 69
rect 111 63 114 66
rect 139 63 142 66
rect 175 63 178 66
rect 187 23 189 63
rect 102 19 105 23
rect 102 14 103 19
rect 102 11 105 14
rect 111 11 114 23
rect 137 19 140 23
rect 157 19 160 23
rect 130 16 140 19
rect 148 16 160 19
rect 130 11 133 16
rect 148 11 151 16
rect 175 11 178 23
rect 200 20 203 23
rect 200 15 208 20
rect 200 11 203 15
rect 218 11 221 23
rect 187 -9 189 11
rect 148 -12 151 -9
rect 148 -15 167 -12
rect 94 -18 99 -17
rect 218 -18 221 -9
rect 90 -25 99 -18
rect 140 -23 142 -18
rect 147 -23 149 -18
rect 140 -25 149 -23
rect 212 -25 221 -18
<< pdm12contact >>
rect 91 23 96 63
rect 118 23 124 63
rect 146 23 151 63
rect 164 23 169 63
rect 189 23 194 63
rect 207 23 212 63
<< psm12contact >>
rect 182 -9 187 11
<< ndm12contact >>
rect 91 -9 96 11
rect 118 -9 124 11
rect 137 -9 142 11
rect 164 -9 169 11
rect 189 -9 194 11
rect 207 -9 212 11
<< nsm12contact >>
rect 182 23 187 63
<< metal2 >>
rect 96 23 118 63
rect 124 23 146 63
rect 151 23 164 63
rect 169 23 182 63
rect 187 23 189 63
rect 194 23 207 63
rect 212 23 221 63
rect 96 -9 118 11
rect 124 -9 137 11
rect 142 -9 164 11
rect 169 -9 182 11
rect 187 -9 189 11
rect 194 -9 207 11
rect 212 -9 221 11
<< labels >>
rlabel metal1 140 -25 149 -18 5 out
rlabel metal1 212 -25 221 -18 5 in
rlabel metal1 189 71 197 77 1 inout
rlabel metal2 109 23 221 63 1 Vdd
rlabel metal2 109 -9 221 11 1 GND
rlabel metal1 90 -25 99 -18 5 oe
rlabel metal1 91 72 99 77 1 oe
<< end >>
