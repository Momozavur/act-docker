magic
tech scmos
timestamp 1764893287
<< error_s >>
rect 97 132 102 133
rect 25 128 30 129
rect 90 16 108 17
rect 90 12 91 16
rect 97 12 103 13
rect 106 12 108 13
rect 25 8 31 9
rect 34 8 36 9
rect 93 -2 99 -1
rect 21 -6 27 -5
rect 97 -25 102 -24
rect 25 -29 30 -28
<< polysilicon >>
rect 120 1202 131 1204
rect 120 1192 131 1194
rect 120 1182 131 1184
rect 120 1171 131 1173
rect 1106 1098 1107 1099
rect 1106 1096 1108 1098
rect 87 1090 89 1094
rect 282 1091 285 1092
rect 1106 941 1107 942
rect 1106 939 1108 941
rect 87 933 89 937
rect 282 934 287 935
rect 1106 784 1107 785
rect 1106 782 1108 784
rect 87 776 89 780
rect 282 777 287 778
rect 1106 627 1107 628
rect 1106 625 1108 627
rect 87 619 89 623
rect 282 620 287 621
rect 1106 470 1107 471
rect 1106 468 1108 470
rect 87 462 89 466
rect 282 463 287 464
rect 1106 313 1107 314
rect 1106 311 1108 313
rect 87 305 89 309
rect 282 306 287 307
rect 1106 156 1107 157
rect 1106 154 1108 156
rect 87 148 89 152
rect 282 149 287 150
rect 1106 -1 1107 0
rect 1106 -3 1108 -1
rect 87 -9 89 -5
rect 282 -8 287 -7
<< polycontact >>
rect 586 1216 591 1221
rect 654 1165 659 1170
rect 1035 1097 1040 1102
rect 12 1087 17 1092
rect 82 1087 87 1092
rect 282 1086 287 1091
rect 519 1087 524 1092
rect 654 1008 659 1013
rect 1035 940 1040 945
rect 12 930 17 935
rect 82 930 87 935
rect 282 929 287 934
rect 519 930 524 935
rect 654 851 659 856
rect 1035 783 1040 788
rect 12 773 17 778
rect 82 773 87 778
rect 282 772 287 777
rect 519 773 524 778
rect 654 694 659 699
rect 1035 626 1040 631
rect 12 616 17 621
rect 82 616 87 621
rect 282 615 287 620
rect 519 616 524 621
rect 654 537 659 542
rect 1035 469 1040 474
rect 12 459 17 464
rect 82 459 87 464
rect 282 458 287 463
rect 519 459 524 464
rect 654 380 659 385
rect 1035 312 1040 317
rect 12 302 17 307
rect 82 302 87 307
rect 282 301 287 306
rect 519 302 524 307
rect 654 223 659 228
rect 1035 155 1040 160
rect 12 145 17 150
rect 82 145 87 150
rect 282 144 287 149
rect 519 145 524 150
rect 654 66 659 71
rect 1035 -2 1040 3
rect 12 -12 17 -7
rect 82 -12 87 -7
rect 282 -13 287 -8
rect 519 -11 524 -6
<< metal1 >>
rect 126 1155 134 1159
rect 122 1154 134 1155
rect 67 1138 72 1154
rect 835 1143 839 1148
rect 937 1143 941 1148
rect 67 1133 116 1138
rect 151 1137 155 1142
rect 1034 1097 1035 1102
rect 74 1084 77 1089
rect 82 1084 87 1087
rect 151 1086 155 1091
rect 344 1084 346 1089
rect 518 1087 519 1092
rect 828 1090 830 1095
rect 351 1063 352 1068
rect 518 1063 523 1087
rect 583 1084 585 1089
rect 1034 1086 1039 1097
rect 1099 1094 1101 1099
rect 929 1081 932 1086
rect 1031 1081 1034 1086
rect 929 1072 932 1077
rect 1031 1072 1034 1077
rect 835 986 839 991
rect 937 986 941 991
rect 151 980 155 985
rect 1034 940 1035 945
rect 74 927 77 932
rect 82 927 87 930
rect 151 929 155 934
rect 344 927 346 932
rect 518 930 519 935
rect 828 933 830 938
rect 351 906 352 911
rect 518 906 523 930
rect 583 927 585 932
rect 1034 929 1039 940
rect 1099 937 1101 942
rect 929 924 932 929
rect 1031 924 1034 929
rect 929 915 932 920
rect 1031 915 1034 920
rect 835 829 839 834
rect 937 829 941 834
rect 151 823 155 828
rect 1034 783 1035 788
rect 74 770 77 775
rect 82 770 87 773
rect 151 772 155 777
rect 344 770 346 775
rect 518 773 519 778
rect 828 776 830 781
rect 351 749 352 754
rect 518 749 523 773
rect 583 770 585 775
rect 1034 772 1039 783
rect 1099 780 1101 785
rect 929 767 932 772
rect 1031 767 1034 772
rect 929 758 932 763
rect 1031 758 1034 763
rect 835 672 839 677
rect 937 672 941 677
rect 151 666 155 671
rect 1034 626 1035 631
rect 74 613 77 618
rect 82 613 87 616
rect 151 615 155 620
rect 344 613 346 618
rect 518 616 519 621
rect 828 619 830 624
rect 351 592 352 597
rect 518 592 523 616
rect 583 613 585 618
rect 1034 615 1039 626
rect 1099 623 1101 628
rect 929 610 932 615
rect 1031 610 1034 615
rect 929 601 932 606
rect 1031 601 1034 606
rect 835 515 839 520
rect 937 515 941 520
rect 151 509 155 514
rect 1034 469 1035 474
rect 74 456 77 461
rect 82 456 87 459
rect 151 458 155 463
rect 344 456 346 461
rect 518 459 519 464
rect 828 462 830 467
rect 351 435 352 440
rect 518 435 523 459
rect 583 456 585 461
rect 1034 458 1039 469
rect 1099 466 1101 471
rect 929 453 932 458
rect 1031 453 1034 458
rect 929 444 932 449
rect 1031 444 1034 449
rect 835 358 839 363
rect 937 358 941 363
rect 151 352 155 357
rect 1034 312 1035 317
rect 74 299 77 304
rect 82 299 87 302
rect 151 301 155 306
rect 344 299 346 304
rect 518 302 519 307
rect 828 305 830 310
rect 351 278 352 283
rect 518 278 523 302
rect 583 299 585 304
rect 1034 301 1039 312
rect 1099 309 1101 314
rect 929 296 932 301
rect 1031 296 1034 301
rect 929 287 932 292
rect 1031 287 1034 292
rect 835 201 839 206
rect 937 201 941 206
rect 151 195 155 200
rect 1034 155 1035 160
rect 74 142 77 147
rect 82 142 87 145
rect 151 144 155 149
rect 344 142 346 147
rect 518 145 519 150
rect 828 148 830 153
rect 351 121 352 126
rect 518 121 523 145
rect 583 142 585 147
rect 1034 144 1039 155
rect 1099 152 1101 157
rect 929 139 932 144
rect 1031 139 1034 144
rect 929 130 932 135
rect 1031 130 1034 135
rect 835 44 839 49
rect 937 44 941 49
rect 151 38 155 43
rect 1034 -2 1035 3
rect 74 -15 77 -10
rect 82 -15 87 -12
rect 151 -13 155 -8
rect 344 -15 346 -10
rect 518 -11 519 -6
rect 828 -9 830 -4
rect 351 -36 352 -31
rect 518 -35 523 -11
rect 583 -15 585 -10
rect 1034 -13 1039 -2
rect 1099 -5 1101 0
rect 929 -18 932 -13
rect 1031 -18 1034 -13
rect 929 -27 932 -22
rect 1031 -27 1034 -22
rect 735 -36 740 -31
<< m2contact >>
rect 932 1143 937 1148
rect 146 1137 151 1142
rect 77 1084 82 1089
rect 346 1084 351 1089
rect 346 1063 351 1068
rect 585 1084 590 1089
rect 1034 1081 1039 1086
rect 932 1072 937 1077
rect 1034 1072 1039 1077
rect 756 1040 761 1058
rect 662 1011 667 1029
rect 932 986 937 991
rect 146 980 151 985
rect 77 927 82 932
rect 346 927 351 932
rect 346 906 351 911
rect 585 927 590 932
rect 1034 924 1039 929
rect 932 915 937 920
rect 1034 915 1039 920
rect 932 829 937 834
rect 146 823 151 828
rect 77 770 82 775
rect 346 770 351 775
rect 346 749 351 754
rect 585 770 590 775
rect 1034 767 1039 772
rect 932 758 937 763
rect 1034 758 1039 763
rect 932 672 937 677
rect 146 666 151 671
rect 77 613 82 618
rect 346 613 351 618
rect 346 592 351 597
rect 585 613 590 618
rect 1034 610 1039 615
rect 932 601 937 606
rect 1034 601 1039 606
rect 932 515 937 520
rect 146 509 151 514
rect 77 456 82 461
rect 346 456 351 461
rect 346 435 351 440
rect 585 456 590 461
rect 1034 453 1039 458
rect 932 444 937 449
rect 1034 444 1039 449
rect 932 358 937 363
rect 146 352 151 357
rect 77 299 82 304
rect 346 299 351 304
rect 346 278 351 283
rect 585 299 590 304
rect 1034 296 1039 301
rect 932 287 937 292
rect 1034 287 1039 292
rect 932 201 937 206
rect 146 195 151 200
rect 77 142 82 147
rect 346 142 351 147
rect 346 121 351 126
rect 585 142 590 147
rect 1034 139 1039 144
rect 932 130 937 135
rect 1034 130 1039 135
rect 932 44 937 49
rect 146 38 151 43
rect 77 -15 82 -10
rect 346 -15 351 -10
rect 346 -36 351 -31
rect 585 -15 590 -10
rect 1034 -18 1039 -13
rect 932 -27 937 -22
rect 1034 -27 1039 -22
<< pm12contact >>
rect 131 1202 136 1207
rect 131 1191 136 1196
rect 131 1180 136 1185
rect 131 1168 136 1173
rect 602 1097 607 1102
rect 764 1094 769 1099
rect 1101 1094 1106 1099
rect 602 940 607 945
rect 764 937 769 942
rect 1101 937 1106 942
rect 602 783 607 788
rect 764 780 769 785
rect 1101 780 1106 785
rect 602 626 607 631
rect 764 623 769 628
rect 1101 623 1106 628
rect 602 469 607 474
rect 764 466 769 471
rect 1101 466 1106 471
rect 602 312 607 317
rect 764 309 769 314
rect 1101 309 1106 314
rect 602 155 607 160
rect 764 152 769 157
rect 1101 152 1106 157
rect 602 -2 607 3
rect 764 -5 769 0
rect 1101 -5 1106 0
<< metal2 >>
rect 839 1175 844 1221
rect 941 1175 946 1221
rect 759 -5 764 0
<< m3contact >>
rect 136 1168 141 1173
<< m123contact >>
rect 1105 1181 1110 1186
rect 649 1165 654 1170
rect 1097 1161 1102 1166
rect 1132 1161 1137 1166
rect 32 1154 37 1159
rect 134 1154 139 1159
rect 830 1143 835 1148
rect 116 1133 121 1138
rect 1124 1141 1129 1146
rect 146 1086 151 1091
rect 830 1090 835 1095
rect 932 1081 937 1086
rect 649 1008 654 1013
rect 830 986 835 991
rect 146 929 151 934
rect 830 933 835 938
rect 932 924 937 929
rect 649 851 654 856
rect 830 829 835 834
rect 146 772 151 777
rect 830 776 835 781
rect 932 767 937 772
rect 649 694 654 699
rect 830 672 835 677
rect 146 615 151 620
rect 830 619 835 624
rect 932 610 937 615
rect 649 537 654 542
rect 830 515 835 520
rect 146 458 151 463
rect 830 462 835 467
rect 932 453 937 458
rect 649 380 654 385
rect 830 358 835 363
rect 146 301 151 306
rect 830 305 835 310
rect 932 296 937 301
rect 649 223 654 228
rect 830 201 835 206
rect 146 144 151 149
rect 830 148 835 153
rect 932 139 937 144
rect 649 66 654 71
rect 830 44 835 49
rect 146 -13 151 -8
rect 830 -9 835 -4
rect 932 -18 937 -13
<< metal3 >>
rect 67 1173 72 1221
rect 155 1188 166 1221
rect 188 1188 199 1221
rect 222 1188 233 1221
rect 255 1188 266 1221
rect 337 1207 342 1221
rect 67 1168 136 1173
rect 30 1154 32 1159
rect 30 1058 35 1154
rect 67 1115 72 1168
rect 116 1118 121 1133
rect 134 1029 139 1154
rect 337 1115 342 1202
rect 439 1175 444 1221
rect 490 1175 495 1221
rect 556 1196 561 1221
rect 556 1185 561 1191
rect 821 1185 826 1221
rect 556 1180 581 1185
rect 576 1115 581 1180
rect 649 1134 654 1165
rect 146 1073 151 1086
rect 649 1073 654 1129
rect 821 1121 826 1180
rect 850 1175 855 1221
rect 923 1175 928 1221
rect 952 1175 957 1221
rect 1025 1175 1030 1221
rect 830 1095 835 1138
rect 932 1091 937 1129
rect 1092 1125 1097 1221
rect 1110 1126 1115 1186
rect 1137 1161 1141 1166
rect 1122 1141 1124 1146
rect 1122 1126 1127 1141
rect 1136 1126 1141 1161
rect 649 977 654 1008
rect 146 916 151 929
rect 649 916 654 972
rect 830 938 835 981
rect 932 934 937 972
rect 649 820 654 851
rect 146 759 151 772
rect 649 759 654 815
rect 830 781 835 824
rect 932 777 937 815
rect 649 663 654 694
rect 146 602 151 615
rect 649 602 654 658
rect 830 624 835 667
rect 932 620 937 658
rect 649 506 654 537
rect 146 445 151 458
rect 649 445 654 501
rect 830 467 835 510
rect 932 463 937 501
rect 649 349 654 380
rect 146 288 151 301
rect 649 288 654 344
rect 830 310 835 353
rect 932 306 937 344
rect 649 192 654 223
rect 146 131 151 144
rect 649 131 654 187
rect 830 153 835 196
rect 932 149 937 187
rect 649 35 654 66
rect 146 -26 151 -13
rect 649 -26 654 30
rect 830 -4 835 39
rect 932 -8 937 30
<< m234contact >>
rect 136 1202 141 1207
rect 136 1191 141 1196
rect 136 1180 141 1185
rect 77 1079 82 1084
rect 146 1142 151 1147
rect 607 1097 612 1102
rect 346 1079 351 1084
rect 585 1079 590 1084
rect 932 1138 937 1143
rect 932 1129 937 1134
rect 1034 1086 1039 1091
rect 1101 1089 1106 1094
rect 346 1068 351 1073
rect 932 1067 937 1072
rect 1034 1067 1039 1072
rect 761 1040 766 1058
rect 667 1011 672 1029
rect 146 985 151 990
rect 607 940 612 945
rect 77 922 82 927
rect 346 922 351 927
rect 585 922 590 927
rect 932 981 937 986
rect 932 972 937 977
rect 1034 929 1039 934
rect 1101 932 1106 937
rect 346 911 351 916
rect 932 910 937 915
rect 1034 910 1039 915
rect 146 828 151 833
rect 607 783 612 788
rect 77 765 82 770
rect 346 765 351 770
rect 585 765 590 770
rect 932 824 937 829
rect 932 815 937 820
rect 1034 772 1039 777
rect 1101 775 1106 780
rect 346 754 351 759
rect 932 753 937 758
rect 1034 753 1039 758
rect 146 671 151 676
rect 607 626 612 631
rect 77 608 82 613
rect 346 608 351 613
rect 585 608 590 613
rect 932 667 937 672
rect 932 658 937 663
rect 1034 615 1039 620
rect 1101 618 1106 623
rect 346 597 351 602
rect 932 596 937 601
rect 1034 596 1039 601
rect 146 514 151 519
rect 607 469 612 474
rect 77 451 82 456
rect 346 451 351 456
rect 585 451 590 456
rect 932 510 937 515
rect 932 501 937 506
rect 1034 458 1039 463
rect 1101 461 1106 466
rect 346 440 351 445
rect 932 439 937 444
rect 1034 439 1039 444
rect 146 357 151 362
rect 607 312 612 317
rect 77 294 82 299
rect 346 294 351 299
rect 585 294 590 299
rect 932 353 937 358
rect 932 344 937 349
rect 1034 301 1039 306
rect 1101 304 1106 309
rect 346 283 351 288
rect 932 282 937 287
rect 1034 282 1039 287
rect 146 200 151 205
rect 607 155 612 160
rect 77 137 82 142
rect 346 137 351 142
rect 585 137 590 142
rect 932 196 937 201
rect 932 187 937 192
rect 1034 144 1039 149
rect 1101 147 1106 152
rect 346 126 351 131
rect 932 125 937 130
rect 1034 125 1039 130
rect 146 43 151 48
rect 607 -2 612 3
rect 77 -20 82 -15
rect 346 -20 351 -15
rect 585 -20 590 -15
rect 932 39 937 44
rect 932 30 937 35
rect 1034 -13 1039 -8
rect 1101 -10 1106 -5
rect 346 -31 351 -26
rect 932 -32 937 -27
rect 1034 -32 1039 -27
<< m4contact >>
rect 337 1202 342 1207
rect 30 1040 35 1058
rect 102 1040 107 1058
rect 556 1191 561 1196
rect 821 1180 826 1185
rect 649 1129 654 1134
rect 830 1138 835 1143
rect 830 1085 835 1090
rect 932 1086 937 1091
rect 146 1068 151 1073
rect 649 1068 654 1073
rect 205 1040 216 1058
rect 300 1039 305 1058
rect 408 1040 413 1059
rect 539 1039 544 1058
rect 784 1040 789 1058
rect 877 1040 882 1058
rect 979 1040 984 1058
rect 1055 1040 1060 1058
rect 1122 1040 1127 1058
rect 18 1011 23 1029
rect 90 1011 95 1029
rect 134 1011 139 1029
rect 270 1011 281 1029
rect 288 1011 293 1029
rect 419 1010 424 1029
rect 527 1011 532 1029
rect 772 1012 777 1030
rect 859 1011 864 1029
rect 961 1011 966 1029
rect 1043 1011 1048 1029
rect 1110 1011 1115 1029
rect 649 972 654 977
rect 830 981 835 986
rect 830 928 835 933
rect 932 929 937 934
rect 146 911 151 916
rect 649 911 654 916
rect 649 815 654 820
rect 830 824 835 829
rect 830 771 835 776
rect 932 772 937 777
rect 146 754 151 759
rect 649 754 654 759
rect 649 658 654 663
rect 830 667 835 672
rect 830 614 835 619
rect 932 615 937 620
rect 146 597 151 602
rect 649 597 654 602
rect 649 501 654 506
rect 830 510 835 515
rect 830 457 835 462
rect 932 458 937 463
rect 146 440 151 445
rect 649 440 654 445
rect 649 344 654 349
rect 830 353 835 358
rect 830 300 835 305
rect 932 301 937 306
rect 146 283 151 288
rect 649 283 654 288
rect 649 187 654 192
rect 830 196 835 201
rect 830 143 835 148
rect 932 144 937 149
rect 146 126 151 131
rect 649 126 654 131
rect 649 30 654 35
rect 830 39 835 44
rect 830 -14 835 -9
rect 932 -13 937 -8
rect 146 -31 151 -26
rect 649 -31 654 -26
<< metal4 >>
rect 141 1202 337 1207
rect 141 1191 556 1196
rect 141 1180 821 1185
rect 131 1168 136 1173
rect 151 1142 608 1147
rect 602 1097 607 1142
rect 835 1138 932 1143
rect 654 1129 932 1134
rect 612 1097 897 1102
rect 830 1084 835 1085
rect 82 1079 346 1084
rect 351 1079 585 1084
rect 590 1079 835 1084
rect 151 1068 346 1073
rect 351 1068 649 1073
rect 892 1072 897 1097
rect 937 1086 1034 1091
rect 1106 1089 1166 1094
rect 892 1067 932 1072
rect 937 1067 1034 1072
rect 35 1040 102 1058
rect 107 1040 205 1058
rect 216 1040 300 1058
rect 305 1040 408 1058
rect 413 1040 539 1058
rect 544 1040 761 1058
rect 766 1040 784 1058
rect 789 1040 877 1058
rect 882 1040 979 1058
rect 984 1040 1055 1058
rect 1060 1040 1122 1058
rect 23 1011 90 1029
rect 95 1011 134 1029
rect 139 1011 270 1029
rect 281 1011 288 1029
rect 293 1011 419 1029
rect 424 1011 527 1029
rect 532 1011 667 1029
rect 672 1012 772 1029
rect 777 1012 859 1029
rect 672 1011 859 1012
rect 864 1011 961 1029
rect 966 1011 1043 1029
rect 1048 1011 1110 1029
rect 151 985 608 990
rect 602 940 607 985
rect 835 981 932 986
rect 654 972 932 977
rect 612 940 897 945
rect 830 927 835 928
rect 82 922 346 927
rect 351 922 585 927
rect 590 922 835 927
rect 151 911 346 916
rect 351 911 649 916
rect 892 915 897 940
rect 937 929 1034 934
rect 1106 932 1166 937
rect 892 910 932 915
rect 937 910 1034 915
rect 151 828 608 833
rect 602 783 607 828
rect 835 824 932 829
rect 654 815 932 820
rect 612 783 897 788
rect 830 770 835 771
rect 82 765 346 770
rect 351 765 585 770
rect 590 765 835 770
rect 151 754 346 759
rect 351 754 649 759
rect 892 758 897 783
rect 937 772 1034 777
rect 1106 775 1166 780
rect 892 753 932 758
rect 937 753 1034 758
rect 151 671 608 676
rect 602 626 607 671
rect 835 667 932 672
rect 654 658 932 663
rect 612 626 897 631
rect 830 613 835 614
rect 82 608 346 613
rect 351 608 585 613
rect 590 608 835 613
rect 151 597 346 602
rect 351 597 649 602
rect 892 601 897 626
rect 937 615 1034 620
rect 1106 618 1166 623
rect 892 596 932 601
rect 937 596 1034 601
rect 151 514 608 519
rect 602 469 607 514
rect 835 510 932 515
rect 654 501 932 506
rect 612 469 897 474
rect 830 456 835 457
rect 82 451 346 456
rect 351 451 585 456
rect 590 451 835 456
rect 151 440 346 445
rect 351 440 649 445
rect 892 444 897 469
rect 937 458 1034 463
rect 1106 461 1166 466
rect 892 439 932 444
rect 937 439 1034 444
rect 151 357 608 362
rect 602 312 607 357
rect 835 353 932 358
rect 654 344 932 349
rect 612 312 897 317
rect 830 299 835 300
rect 82 294 346 299
rect 351 294 585 299
rect 590 294 835 299
rect 151 283 346 288
rect 351 283 649 288
rect 892 287 897 312
rect 937 301 1034 306
rect 1106 304 1166 309
rect 892 282 932 287
rect 937 282 1034 287
rect 151 200 608 205
rect 602 155 607 200
rect 835 196 932 201
rect 654 187 932 192
rect 612 155 897 160
rect 830 142 835 143
rect 82 137 346 142
rect 351 137 585 142
rect 590 137 835 142
rect 151 126 346 131
rect 351 126 649 131
rect 892 130 897 155
rect 937 144 1034 149
rect 1106 147 1166 152
rect 892 125 932 130
rect 937 125 1034 130
rect 151 43 608 48
rect 602 -2 607 43
rect 835 39 932 44
rect 654 30 932 35
rect 612 -2 897 3
rect 830 -15 835 -14
rect 82 -20 346 -15
rect 351 -20 585 -15
rect 590 -20 835 -15
rect 151 -31 346 -26
rect 351 -31 649 -26
rect 892 -27 897 -2
rect 937 -13 1034 -8
rect 1106 -10 1166 -5
rect 892 -32 932 -27
rect 937 -32 1034 -27
use 4nor  4nor_0
timestamp 1761285742
transform 0 1 53 -1 0 1289
box 68 -24 135 80
use staticizer  staticizer_0
timestamp 1761284585
transform 1 0 26 0 1 1063
box 61 -1099 120 61
use fblock  fblock_0
timestamp 1761104028
transform 1 0 161 0 1 1041
box -6 -1077 124 175
use latch  latch_0
timestamp 1761111742
transform 1 0 407 0 1 -120
box -392 84 -333 1235
use latch  latch_1
timestamp 1761111742
transform 1 0 677 0 1 -120
box -392 84 -333 1235
use shift  shift_0
timestamp 1761107410
transform 1 0 442 0 1 325
box -90 -361 79 853
use latch  latch_2
timestamp 1761111742
transform 1 0 916 0 1 -120
box -392 84 -333 1235
use addsub  addsub_0
timestamp 1761186134
transform 1 0 598 0 1 4
box -7 -40 166 1226
use reg  reg_0
timestamp 1761104463
transform 1 0 853 0 1 369
box -14 -399 76 806
use latch  latch_3
timestamp 1761111742
transform 1 0 1161 0 1 -114
box -392 84 -333 1235
use reg  reg_1
timestamp 1761104463
transform 1 0 955 0 1 369
box -14 -399 76 806
use latch  latch_4
timestamp 1761111742
transform 1 0 1432 0 1 -110
box -392 84 -333 1235
use staticizer  staticizer_1
timestamp 1761284585
transform 1 0 1046 0 1 1065
box 61 -1099 120 61
use inv  inv_0
timestamp 1758863638
transform 1 0 1112 0 1 1150
box -10 -12 20 39
<< labels >>
rlabel metal3 1136 1151 1141 1155 1 stat2_en
rlabel metal4 161 -31 166 -26 1 rx7
rlabel metal4 161 126 166 131 1 rx6
rlabel metal4 161 283 166 288 1 rx5
rlabel metal4 161 440 166 445 1 rx4
rlabel metal4 161 597 166 602 1 rx3
rlabel metal4 161 754 166 759 1 rx2
rlabel metal4 161 911 166 916 1 rx1
rlabel metal4 161 1068 166 1073 1 rx0
rlabel metal4 165 985 170 990 1 ry1
rlabel metal4 165 43 170 48 1 ry7
rlabel metal4 165 200 170 205 1 ry6
rlabel metal4 165 357 170 362 1 ry5
rlabel metal4 165 514 170 519 1 ry4
rlabel metal4 165 671 170 676 1 ry3
rlabel metal4 165 828 170 833 1 ry2
rlabel metal4 165 1142 170 1147 1 ry0
rlabel metal4 97 -20 102 -15 1 wz7
rlabel metal4 97 137 102 142 1 wz6
rlabel metal4 97 294 102 299 1 wz5
rlabel metal4 97 451 102 456 1 wz4
rlabel metal4 97 608 102 613 1 wz3
rlabel metal4 97 765 102 770 1 wz2
rlabel metal4 97 922 102 927 1 wz1
rlabel metal4 97 1079 102 1084 1 wz0
rlabel metal4 1161 1089 1166 1094 7 out0
rlabel metal4 1161 932 1166 937 7 out1
rlabel metal4 1161 775 1166 780 7 out2
rlabel metal4 1161 618 1166 623 7 out3
rlabel metal4 1161 461 1166 466 7 out4
rlabel metal4 1161 304 1166 309 7 out5
rlabel metal4 1161 147 1166 152 7 out6
rlabel metal4 1161 -10 1166 -5 7 out7
rlabel m4contact 18 1011 23 1029 1 Vdd!
rlabel m4contact 30 1040 35 1058 1 GND!
rlabel polycontact 12 -12 17 -7 3 in7
rlabel polycontact 12 145 17 150 3 in6
rlabel polycontact 12 302 17 307 3 in5
rlabel polycontact 12 459 17 464 3 in4
rlabel polycontact 12 616 17 621 3 in3
rlabel polycontact 12 773 17 778 3 in2
rlabel polycontact 12 930 17 935 3 in1
rlabel polycontact 12 1087 17 1092 3 in0
rlabel metal3 1092 1216 1097 1221 1 rd
rlabel metal3 821 1216 826 1221 1 ras
rlabel metal3 556 1216 561 1221 1 ros
rlabel metal3 337 1216 342 1221 1 rfb
rlabel metal1 735 -36 740 -31 1 as_cout
rlabel polycontact 586 1216 591 1221 1 as_cin
rlabel metal3 490 1216 495 1221 1 os_s
rlabel metal3 439 1216 444 1221 1 os_u
rlabel metal3 255 1216 266 1221 1 fb_g0
rlabel metal3 222 1216 233 1221 1 fb_g1
rlabel metal3 188 1216 199 1221 1 fb_g2
rlabel metal3 155 1216 166 1221 1 fb_g3
rlabel metal3 1025 1216 1030 1221 1 reg1_w
rlabel metal3 952 1216 957 1221 1 reg1_r1
rlabel metal2 941 1216 946 1221 1 reg1_r0
rlabel metal3 923 1216 928 1221 1 reg0_w
rlabel metal3 850 1216 855 1221 1 reg0_r1
rlabel metal2 839 1216 844 1221 1 reg0_r0
rlabel metal3 67 1216 72 1221 1 ld
<< end >>
