magic
tech scmos
timestamp 1765780088
<< metal5 >>
rect -108 90 -88 94
rect -108 82 -104 90
rect -92 82 -88 90
rect -108 78 -88 82
rect -84 90 -62 94
rect -84 82 -80 90
rect -66 82 -62 90
rect -84 78 -62 82
rect -58 90 -36 94
rect -58 82 -54 90
rect -40 82 -36 90
rect -58 78 -36 82
rect -108 64 -104 78
rect -84 74 -72 78
rect -84 64 -80 74
rect -76 70 -68 74
rect -72 66 -64 70
rect -68 64 -64 66
rect -58 64 -54 78
rect -40 64 -36 78
rect -32 90 -18 94
rect -10 90 -6 94
rect 8 90 12 94
rect -32 68 -28 90
rect -22 86 -14 90
rect -10 86 -2 90
rect 4 86 12 90
rect -18 72 -14 86
rect -6 82 8 86
rect -22 68 -14 72
rect -32 64 -18 68
rect -1 64 3 82
rect 16 68 20 94
rect 34 68 38 94
rect 16 64 38 68
rect 42 90 46 94
rect 42 86 50 90
rect 42 82 54 86
rect 42 64 46 82
rect 50 78 56 82
rect 60 78 64 94
rect 52 74 64 78
rect 88 90 106 94
rect 110 90 132 94
rect 88 81 92 90
rect 88 77 106 81
rect 58 70 64 74
rect 60 64 64 70
rect 102 68 106 77
rect 88 64 106 68
rect 110 68 114 90
rect 128 68 132 90
rect 110 64 132 68
rect 136 68 140 94
rect 158 90 176 94
rect 182 90 196 94
rect 158 82 162 90
rect 172 82 176 90
rect 158 78 176 82
rect 136 64 154 68
rect 158 64 162 78
rect 172 64 176 78
rect 188 68 192 90
rect 182 64 196 68
rect -128 36 -112 40
rect -128 28 -124 36
rect -116 28 -112 36
rect -128 24 -112 28
rect -128 10 -124 24
rect -116 10 -112 24
rect -108 36 -104 40
rect -108 32 -100 36
rect -108 28 -96 32
rect -108 10 -104 28
rect -100 27 -96 28
rect -100 23 -94 27
rect -98 22 -94 23
rect -90 22 -86 40
rect -82 36 -60 40
rect -56 36 -40 40
rect -98 18 -86 22
rect -94 14 -86 18
rect -90 10 -86 14
rect -73 10 -69 36
rect -56 14 -52 36
rect -44 14 -40 36
rect -56 10 -40 14
rect -36 36 -32 40
rect -36 32 -28 36
rect -36 28 -24 32
rect -36 10 -32 28
rect -28 27 -24 28
rect -28 23 -22 27
rect -26 22 -22 23
rect -18 22 -14 40
rect -26 18 -14 22
rect -22 14 -14 18
rect -18 10 -14 14
rect 10 36 14 40
rect 26 36 30 40
rect 10 32 18 36
rect 22 32 30 36
rect 10 28 30 32
rect 10 10 14 28
rect 18 24 22 28
rect 26 10 30 28
rect 34 36 56 40
rect 34 27 38 36
rect 34 23 56 27
rect 34 14 38 23
rect 60 14 64 40
rect 82 36 86 40
rect 82 32 90 36
rect 82 28 94 32
rect 34 10 56 14
rect 60 10 78 14
rect 82 10 86 28
rect 90 26 95 28
rect 90 24 96 26
rect 91 22 96 24
rect 100 22 104 40
rect 108 36 112 40
rect 124 36 128 40
rect 108 32 116 36
rect 120 32 128 36
rect 132 36 150 40
rect 112 28 124 32
rect 92 18 104 22
rect 96 14 104 18
rect 100 10 104 14
rect 116 10 120 28
rect 132 14 136 36
rect 154 28 158 40
rect 168 28 172 40
rect 154 24 172 28
rect 132 10 150 14
rect 154 10 158 24
rect 168 10 172 24
rect 176 14 180 40
rect 194 14 198 40
rect 176 10 198 14
rect 202 27 206 40
rect 218 35 222 40
rect 214 31 222 35
rect 210 27 218 31
rect 202 23 214 27
rect 202 10 206 23
rect 210 19 218 23
rect 214 15 222 19
rect 218 10 222 15
rect -103 -18 -99 -14
rect -87 -18 -83 -14
rect -103 -22 -95 -18
rect -91 -22 -83 -18
rect -103 -26 -83 -22
rect -103 -44 -99 -26
rect -95 -30 -91 -26
rect -87 -44 -83 -26
rect -79 -18 -57 -14
rect -79 -40 -75 -18
rect -61 -40 -57 -18
rect -79 -44 -57 -40
rect -53 -18 -49 -14
rect -37 -18 -33 -14
rect -53 -22 -45 -18
rect -41 -22 -33 -18
rect -53 -26 -33 -22
rect -53 -44 -49 -26
rect -45 -30 -41 -26
rect -37 -44 -33 -26
rect -29 -18 -11 -14
rect -29 -40 -25 -18
rect -7 -26 -3 -14
rect 7 -26 11 -14
rect 15 -18 29 -14
rect -7 -30 11 -26
rect -29 -44 -11 -40
rect -7 -44 -3 -30
rect 7 -44 11 -30
rect 21 -40 25 -18
rect 33 -40 37 -14
rect 75 -26 79 -14
rect 93 -18 97 -14
rect 89 -22 97 -18
rect 101 -18 123 -14
rect 85 -26 93 -22
rect 75 -30 89 -26
rect 15 -44 29 -40
rect 33 -44 51 -40
rect 75 -44 79 -30
rect 85 -34 93 -30
rect 89 -38 97 -34
rect 93 -44 97 -38
rect 101 -40 105 -18
rect 119 -40 123 -18
rect 101 -44 123 -40
rect 127 -40 131 -14
rect 149 -18 167 -14
rect 149 -26 153 -18
rect 149 -30 165 -26
rect 149 -40 153 -30
rect 171 -36 175 -14
rect 185 -36 189 -14
rect 171 -40 189 -36
rect 127 -44 145 -40
rect 149 -44 167 -40
rect 175 -44 185 -40
<< end >>
