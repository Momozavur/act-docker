magic
tech scmos
timestamp 1765697223
<< polysilicon >>
rect 175 32 177 41
rect 186 32 188 41
rect 175 -38 177 -29
rect 186 -38 188 -29
rect 175 -108 177 -99
rect 186 -108 188 -99
rect 175 -178 177 -169
rect 186 -178 188 -169
<< polycontact >>
rect 184 41 189 46
rect 184 -29 189 -24
rect 184 -99 189 -94
rect 184 -169 189 -164
<< metal1 >>
rect 114 -94 119 56
rect 114 -164 119 -99
rect 114 -312 119 -169
rect 124 46 129 56
rect 124 -24 129 41
rect 124 -273 129 -29
rect 134 -14 139 56
rect 134 -154 139 -19
rect 134 -263 139 -159
rect 144 51 189 56
rect 144 -84 149 51
rect 184 46 189 51
rect 184 -24 189 -19
rect 144 -89 189 -84
rect 144 -224 149 -89
rect 184 -94 189 -89
rect 184 -164 189 -159
rect 144 -229 173 -224
rect 168 -231 173 -229
rect 186 -234 191 -214
rect 168 -263 173 -254
rect 134 -268 173 -263
rect 124 -278 153 -273
rect 186 -274 191 -255
rect 148 -280 153 -278
rect 166 -279 191 -274
rect 166 -284 171 -279
rect 148 -312 153 -308
rect 114 -317 153 -312
<< m2contact >>
rect 114 -169 119 -164
rect 124 41 129 46
rect 124 -29 129 -24
rect 134 -19 139 -14
rect 134 -159 139 -154
rect 209 33 214 38
rect 199 -9 204 -4
rect 184 -19 189 -14
rect 209 -37 214 -32
rect 199 -79 204 -74
rect 209 -107 214 -102
rect 199 -149 204 -144
rect 184 -159 189 -154
rect 209 -177 214 -172
rect 199 -219 204 -214
rect 144 -248 149 -243
rect 124 -295 129 -290
<< pm12contact >>
rect 114 -99 119 -94
rect 174 41 179 46
rect 174 -29 179 -24
rect 174 -99 179 -94
rect 174 -169 179 -164
<< metal2 >>
rect 129 41 174 46
rect 139 -19 184 -14
rect 129 -29 174 -24
rect 199 -74 204 -9
rect 119 -99 174 -94
rect 199 -144 204 -79
rect 139 -159 184 -154
rect 119 -169 174 -164
rect 199 -214 204 -149
rect 209 -32 214 33
rect 209 -102 214 -37
rect 209 -172 214 -107
rect 209 -243 214 -177
rect 124 -248 144 -243
rect 149 -248 214 -243
rect 124 -290 129 -248
use 2and  2and_0
timestamp 1765690562
transform 1 0 90 0 1 -41
box 68 29 138 82
use 2and  2and_3
timestamp 1765690562
transform 1 0 90 0 1 -251
box 68 29 138 82
use 2and  2and_2
timestamp 1765690562
transform 1 0 90 0 1 -181
box 68 29 138 82
use 2and  2and_1
timestamp 1765690562
transform 1 0 90 0 1 -111
box 68 29 138 82
use inv2  inv2_0
timestamp 1765338958
transform 0 -1 161 1 0 -298
box -10 -13 20 40
use inv2  inv2_1
timestamp 1765338958
transform 0 -1 181 1 0 -251
box -10 -13 20 40
<< end >>
