magic
tech scmos
timestamp 1765416915
use 2mux_nr  2mux_nr_2 /home/user
timestamp 1765248526
transform 0 -1 22 -1 0 -61
box -32 -38 29 27
use 2mux_nr  2mux_nr_0
timestamp 1765248526
transform 0 -1 22 -1 0 0
box -32 -38 29 27
use 2mux_nr  2mux_nr_1
timestamp 1765248526
transform 0 -1 87 -1 0 0
box -32 -38 29 27
use inv  inv_0 /home/user
timestamp 1765001281
transform 1 0 73 0 1 -76
box -10 -13 20 40
use inv  inv_2
timestamp 1765001281
transform 1 0 38 0 1 46
box -10 -13 20 40
use inv  inv_4
timestamp 1765001281
transform 1 0 105 0 1 46
box -10 -13 20 40
use inv  inv_1
timestamp 1765001281
transform 1 0 5 0 1 46
box -10 -13 20 40
use inv  inv_3
timestamp 1765001281
transform 1 0 72 0 1 46
box -10 -13 20 40
<< labels >>
rlabel metal1 0 59 0 59 3 g3
rlabel metal1 32 59 32 59 1 g2
rlabel metal1 66 60 66 60 1 g1
rlabel metal1 101 58 101 58 1 g0
rlabel metal1 91 -43 91 -43 1 f
rlabel metal1 -3 -63 -3 -63 3 a
rlabel metal1 -3 -3 -3 -3 3 b
rlabel metal1 32 38 32 38 1 GND!
rlabel metal1 25 80 25 80 1 Vdd!
<< end >>
