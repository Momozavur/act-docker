magic
tech scmos
timestamp 1765001281
<< nwell >>
rect -10 14 20 40
<< pwell >>
rect -10 -13 20 13
<< ntransistor >>
rect 4 0 6 7
<< ptransistor >>
rect 4 20 6 27
<< ndiffusion >>
rect 1 0 4 7
rect 6 0 9 7
<< pdiffusion >>
rect 1 20 4 27
rect 6 20 9 27
<< ndcontact >>
rect -4 0 1 7
rect 9 0 14 7
<< pdcontact >>
rect -4 20 1 27
rect 9 20 14 27
<< psubstratepcontact >>
rect -2 -10 12 -5
<< nsubstratencontact >>
rect -2 32 12 37
<< polysilicon >>
rect 4 27 6 30
rect 4 16 6 20
rect 4 7 6 11
rect 4 -3 6 0
<< polycontact >>
rect 1 11 6 16
<< metal1 >>
rect -7 32 -2 37
rect 12 32 17 37
rect -4 27 1 32
rect 9 16 14 20
rect -10 11 1 16
rect 9 11 20 16
rect 9 7 14 11
rect -4 -5 1 0
rect -7 -10 -2 -5
rect 12 -10 17 -5
<< labels >>
rlabel metal1 -10 11 -10 16 3 in
rlabel metal1 20 11 20 16 7 out
rlabel metal1 -5 34 -5 34 3 Vdd!
rlabel metal1 -5 -7 -5 -7 3 GND!
<< end >>
