magic
tech scmos
timestamp 1765795763
<< pwell >>
rect 879 3604 884 3620
rect 1229 3604 1234 3620
rect 1489 1638 1494 1643
rect 1234 1616 1235 1625
<< polysilicon >>
rect 1684 3210 1686 3223
rect 1611 3198 1669 3200
rect 1621 3187 1669 3189
rect 1631 3176 1669 3178
rect 1684 3043 1686 3046
rect 1656 2983 1657 2985
rect 1655 2958 1657 2983
rect 1683 2969 1685 2981
rect 1655 2956 1669 2958
rect 1298 1802 1300 1815
rect 1309 1802 1311 1815
<< polycontact >>
rect 1684 3223 1689 3228
rect 1606 3198 1611 3203
rect 1616 3187 1621 3192
rect 1626 3176 1631 3181
rect 1685 3162 1690 3167
rect 1684 3102 1689 3107
rect 1681 3046 1686 3051
rect 1651 2983 1656 2988
rect 1681 2981 1686 2986
rect 1832 1790 1837 1795
rect 2332 1790 2337 1795
<< metal1 >>
rect 75 3403 314 3411
rect 75 3053 283 3062
rect 270 2750 283 3053
rect 301 2781 314 3403
rect 656 3341 665 3597
rect 3309 3353 3587 3490
rect 3309 3348 3310 3353
rect 3348 3348 3587 3353
rect 656 3331 1668 3341
rect 1658 3282 1668 3331
rect 2644 3285 2649 3286
rect 1331 3254 1351 3259
rect 1663 3217 1668 3227
rect 1705 3217 1710 3227
rect 1662 3158 1667 3168
rect 1685 3167 1690 3169
rect 1706 3160 1711 3168
rect 1711 3149 1721 3154
rect 2460 3134 2465 3139
rect 1649 3125 1667 3130
rect 1649 3089 1655 3125
rect 1682 3102 1684 3107
rect 1649 3084 1665 3089
rect 2470 3087 2475 3092
rect 1664 3047 1669 3066
rect 1661 3042 1669 3047
rect 1474 2925 1479 2930
rect 1474 2861 1479 2866
rect 1474 2797 1479 2802
rect 1679 2796 1684 2925
rect 3575 2792 3623 2799
rect 3575 2781 3582 2792
rect 301 2772 360 2781
rect 270 2741 339 2750
rect 75 2703 324 2712
rect 297 2362 306 2363
rect 75 2353 306 2362
rect 75 2003 290 2012
rect 279 1968 290 2003
rect 72 1652 267 1663
rect 255 1562 267 1652
rect 224 1312 235 1314
rect 73 1303 235 1312
rect 74 953 205 962
rect 194 612 205 953
rect 224 612 235 1303
rect 256 689 266 1562
rect 279 1485 288 1968
rect 278 864 288 1485
rect 297 1240 306 2353
rect 296 1170 306 1240
rect 315 1408 324 2703
rect 330 1586 339 2741
rect 315 1216 325 1408
rect 330 1392 340 1586
rect 349 1566 360 2772
rect 3575 2776 3583 2781
rect 1474 2733 1479 2738
rect 2308 2704 2317 2713
rect 455 2695 464 2704
rect 455 2263 464 2686
rect 455 2244 464 2254
rect 569 2677 578 2704
rect 569 2262 578 2668
rect 569 2244 578 2253
rect 683 2659 692 2704
rect 683 2263 692 2650
rect 683 2245 692 2254
rect 797 2641 806 2704
rect 797 2263 806 2632
rect 797 2245 806 2254
rect 911 2623 920 2704
rect 911 2263 920 2614
rect 911 2245 920 2254
rect 1025 2605 1034 2704
rect 1025 2263 1034 2596
rect 1025 2245 1034 2254
rect 1139 2587 1148 2704
rect 1139 2263 1148 2578
rect 1139 2245 1148 2254
rect 1253 2569 1262 2704
rect 2380 2595 2385 2600
rect 3445 2561 3477 2562
rect 1253 2263 1262 2560
rect 2360 2546 2365 2551
rect 3258 2516 3477 2561
rect 1253 2245 1262 2254
rect 2608 2257 2617 2266
rect 2608 2248 2660 2257
rect 1253 1758 1258 1784
rect 1805 1769 1814 1774
rect 2305 1769 2316 1774
rect 1253 1753 1278 1758
rect 1273 1634 1278 1753
rect 1286 1727 1291 1762
rect 1805 1729 1810 1769
rect 1805 1724 1816 1729
rect 1835 1725 1840 1732
rect 2305 1729 2310 1769
rect 2609 1737 2618 1764
rect 2305 1724 2316 1729
rect 2335 1722 2340 1737
rect 2609 1732 2640 1737
rect 2651 1732 2660 2248
rect 2611 1729 2616 1732
rect 2653 1728 2658 1732
rect 3130 1535 3135 1540
rect 3254 1535 3259 1540
rect 330 1384 351 1392
rect 333 1383 351 1384
rect 3130 1359 3135 1364
rect 3254 1359 3259 1364
rect 315 1214 353 1216
rect 315 1209 356 1214
rect 315 1207 353 1209
rect 315 1206 325 1207
rect 3130 1183 3135 1188
rect 3254 1183 3259 1188
rect 296 1040 305 1170
rect 296 1038 351 1040
rect 296 1033 356 1038
rect 296 1031 351 1033
rect 3130 1007 3135 1012
rect 3254 1007 3259 1012
rect 278 862 351 864
rect 278 857 356 862
rect 278 855 351 857
rect 3130 831 3135 836
rect 3254 831 3259 836
rect 256 688 348 689
rect 256 686 351 688
rect 256 681 356 686
rect 256 680 351 681
rect 256 679 284 680
rect 342 679 351 680
rect 256 678 266 679
rect 3130 655 3135 660
rect 3254 655 3259 660
rect 68 542 75 555
rect 87 542 93 581
rect 27 536 93 542
rect 194 337 205 603
rect 224 513 235 603
rect 224 512 297 513
rect 224 510 351 512
rect 224 505 356 510
rect 224 503 351 505
rect 224 502 235 503
rect 3130 479 3135 484
rect 3254 479 3259 484
rect 194 336 238 337
rect 194 334 351 336
rect 194 329 356 334
rect 194 327 351 329
rect 194 326 238 327
rect 3130 303 3135 308
rect 3254 303 3259 308
rect 3445 90 3477 2516
rect 3575 2442 3623 2449
rect 3575 2431 3582 2442
rect 3575 2426 3583 2431
rect 3575 2092 3623 2099
rect 3575 2081 3582 2092
rect 3575 2076 3583 2081
rect 3575 1742 3623 1749
rect 3575 1731 3582 1742
rect 3575 1726 3583 1731
rect 3575 1392 3623 1399
rect 3575 1381 3582 1392
rect 3575 1376 3583 1381
rect 3575 1042 3623 1049
rect 3575 1031 3582 1042
rect 3575 1026 3583 1031
rect 3575 692 3623 699
rect 3575 681 3582 692
rect 3575 676 3583 681
rect 3575 342 3623 349
rect 3575 335 3582 342
<< m2contact >>
rect 534 3585 543 3594
rect 75 3475 84 3484
rect 75 3125 84 3134
rect 75 2775 84 2784
rect 884 3585 893 3594
rect 1234 3585 1243 3594
rect 1356 3585 1365 3594
rect 3310 3347 3348 3353
rect 1658 3273 1668 3282
rect 3206 3273 3212 3279
rect 1344 3246 1353 3254
rect 1596 3253 1601 3258
rect 1684 3253 1689 3258
rect 1705 3096 1710 3101
rect 1666 3007 1671 3012
rect 1667 2975 1672 2980
rect 1351 2896 1360 2905
rect 1351 2832 1360 2841
rect 1679 2791 1684 2796
rect 2344 2786 2353 2795
rect 3623 2792 3630 2799
rect 75 2425 84 2434
rect 75 2075 84 2084
rect 75 1725 84 1734
rect 75 1375 84 1384
rect 75 1025 84 1034
rect 87 628 93 634
rect 1351 2768 1360 2777
rect 3566 2726 3575 2735
rect 1351 2704 1360 2713
rect 2317 2704 2326 2713
rect 455 2686 464 2695
rect 569 2668 578 2677
rect 683 2650 692 2659
rect 797 2632 806 2641
rect 911 2614 920 2623
rect 1025 2596 1034 2605
rect 1139 2578 1148 2587
rect 1253 2560 1262 2569
rect 2608 2266 2617 2275
rect 1317 1799 1322 1804
rect 2609 1764 2618 1773
rect 1853 1716 1858 1721
rect 1489 1638 1494 1643
rect 3186 1564 3194 1572
rect 3310 1548 3318 1557
rect 1959 1523 1964 1528
rect 3186 1388 3194 1396
rect 3310 1372 3318 1381
rect 1959 1347 1964 1352
rect 3186 1212 3194 1220
rect 3310 1196 3318 1205
rect 1959 1171 1964 1176
rect 3186 1036 3194 1044
rect 3310 1020 3318 1029
rect 1959 995 1964 1000
rect 3186 860 3194 868
rect 3310 844 3318 853
rect 1959 819 1964 824
rect 3186 684 3194 692
rect 3310 668 3318 677
rect 1959 643 1964 648
rect 20 536 27 542
rect 3186 508 3194 516
rect 3310 492 3318 501
rect 1959 467 1964 472
rect 3186 332 3194 340
rect 3310 316 3318 325
rect 1959 291 1964 296
rect 607 94 616 102
rect 957 94 966 102
rect 1307 94 1316 102
rect 1657 94 1666 102
rect 2007 94 2016 102
rect 2357 94 2366 102
rect 2707 94 2716 102
rect 3057 94 3066 102
rect 3623 2442 3630 2449
rect 3566 2376 3575 2385
rect 3623 2092 3630 2099
rect 3566 2026 3575 2035
rect 3623 1742 3630 1749
rect 3566 1676 3575 1685
rect 3623 1392 3630 1399
rect 3566 1326 3575 1335
rect 3623 1042 3630 1049
rect 3566 976 3575 985
rect 3623 692 3630 699
rect 3566 626 3575 635
rect 3623 342 3630 349
rect 3566 276 3575 285
<< pm12contact >>
rect 1296 1815 1301 1820
rect 1309 1815 1314 1820
<< metal2 >>
rect 525 3585 534 3620
rect 875 3585 884 3620
rect 1225 3585 1234 3620
rect 84 3475 331 3484
rect 84 3125 313 3134
rect 84 2775 296 2784
rect 286 2680 296 2775
rect 286 2659 295 2680
rect 304 2677 313 3125
rect 322 2695 331 3475
rect 1356 3307 1365 3585
rect 1344 3299 1365 3307
rect 3206 3347 3310 3352
rect 3348 3347 3349 3352
rect 3206 3346 3349 3347
rect 340 3259 345 3262
rect 448 3259 453 3262
rect 603 3259 608 3262
rect 749 3259 754 3262
rect 1344 3254 1353 3299
rect 3206 3279 3212 3346
rect 1601 3253 1684 3258
rect 1671 3007 1674 3012
rect 1669 2980 1674 3007
rect 1672 2975 1674 2980
rect 1705 2972 1710 3096
rect 528 2800 533 2803
rect 642 2800 647 2803
rect 756 2799 761 2802
rect 870 2800 875 2803
rect 984 2800 989 2803
rect 1212 2799 1217 2802
rect 1326 2799 1331 2802
rect 1098 2785 1103 2788
rect 322 2686 455 2695
rect 304 2668 569 2677
rect 286 2650 683 2659
rect 258 2632 797 2641
rect 258 2434 267 2632
rect 84 2425 267 2434
rect 276 2614 911 2623
rect 276 2084 285 2614
rect 84 2075 285 2084
rect 294 2596 1025 2605
rect 294 1734 303 2596
rect 84 1725 303 1734
rect 312 2578 1139 2587
rect 312 1725 321 2578
rect 313 1384 321 1725
rect 84 1375 321 1384
rect 330 2560 1253 2569
rect 330 1034 339 2560
rect 2598 2225 2603 2232
rect 1317 1754 1322 1799
rect 1848 1770 1862 1775
rect 2348 1770 2362 1775
rect 2594 1773 2603 2225
rect 1848 1716 1853 1770
rect 2348 1716 2353 1770
rect 2594 1764 2609 1773
rect 2681 1764 2690 2214
rect 2699 2205 2708 2222
rect 2699 1764 2708 2196
rect 2717 2187 2726 2222
rect 2717 1764 2726 2178
rect 2735 2169 2744 2222
rect 2735 1764 2744 2160
rect 2763 2151 2772 2222
rect 2763 1764 2772 2142
rect 2781 2133 2790 2222
rect 2781 1764 2790 2124
rect 2799 2115 2808 2222
rect 2799 1764 2808 2106
rect 2817 2097 2826 2222
rect 2817 1764 2826 2088
rect 2845 2079 2854 2222
rect 2845 1764 2854 2070
rect 2863 2061 2872 2222
rect 2863 1764 2872 2052
rect 2881 2043 2890 2222
rect 2881 1764 2890 2034
rect 2899 2025 2908 2222
rect 2899 1764 2908 2016
rect 2927 2007 2936 2222
rect 2927 1764 2936 1998
rect 2945 1989 2954 2222
rect 2945 1764 2954 1980
rect 2963 1971 2972 2222
rect 2963 1764 2972 1962
rect 2981 1953 2990 2222
rect 2981 1764 2990 1944
rect 3009 1935 3018 2222
rect 3009 1755 3018 1926
rect 3027 1917 3036 2222
rect 3027 1765 3036 1908
rect 3045 1899 3054 2222
rect 2384 1746 3018 1755
rect 3045 1737 3054 1890
rect 3063 1881 3072 2222
rect 3063 1764 3072 1872
rect 3091 1863 3100 2222
rect 3091 1764 3100 1854
rect 3109 1845 3118 2222
rect 3109 1764 3118 1836
rect 3127 1827 3136 2222
rect 3127 1764 3136 1818
rect 3145 1809 3154 2222
rect 3145 1764 3154 1800
rect 3173 1791 3182 2222
rect 3173 1764 3182 1782
rect 3189 1773 3198 2222
rect 3209 1791 3218 2222
rect 3209 1764 3218 1782
rect 3227 1764 3236 2222
rect 3000 1728 3054 1737
rect 3000 1697 3009 1728
rect 2364 1688 3009 1697
rect 715 1612 782 1617
rect 1452 1612 1457 1616
rect 1559 1612 1564 1616
rect 1666 1612 1671 1616
rect 2364 1617 2373 1688
rect 1866 1612 1871 1615
rect 2366 1615 2373 1617
rect 2366 1612 2371 1615
rect 2473 1612 2478 1616
rect 2666 1612 2671 1616
rect 804 1611 864 1612
rect 804 1607 859 1611
rect 2661 1607 2671 1612
rect 3000 1608 3009 1688
rect 84 1025 339 1034
rect 59 697 93 704
rect 87 634 93 697
<< m3contact >>
rect 1582 2967 1587 2972
rect 2681 2214 2690 2223
rect 2699 2196 2708 2205
rect 2717 2178 2726 2187
rect 2735 2160 2744 2169
rect 2763 2142 2772 2151
rect 2781 2124 2790 2133
rect 2799 2106 2808 2115
rect 2817 2088 2826 2097
rect 2845 2070 2854 2079
rect 2863 2052 2872 2061
rect 2881 2034 2890 2043
rect 2899 2016 2908 2025
rect 2927 1998 2936 2007
rect 2945 1980 2954 1989
rect 2963 1962 2972 1971
rect 2981 1944 2990 1953
rect 3009 1926 3018 1935
rect 3027 1908 3036 1917
rect 3045 1890 3054 1899
rect 2375 1746 2384 1755
rect 3063 1872 3072 1881
rect 3091 1854 3100 1863
rect 3109 1836 3118 1845
rect 3127 1818 3136 1827
rect 3145 1800 3154 1809
rect 3173 1782 3182 1791
rect 3189 1764 3198 1773
rect 3209 1782 3218 1791
rect 1559 1616 1564 1621
rect 1666 1616 1671 1621
<< m123contact >>
rect 75 3353 84 3362
rect 75 3003 84 3012
rect 75 2653 84 2662
rect 2591 3285 2597 3291
rect 2644 3286 2649 3291
rect 1714 3128 1719 3133
rect 1738 3128 1743 3133
rect 1717 3107 1722 3112
rect 1663 3089 1668 3094
rect 1651 3075 1656 3080
rect 1646 2983 1651 2988
rect 1705 2967 1710 2972
rect 1663 2948 1668 2953
rect 2367 2883 2376 2892
rect 75 2303 84 2312
rect 75 1953 84 1962
rect 75 1603 84 1612
rect 75 1253 84 1262
rect 455 2254 464 2263
rect 569 2253 578 2262
rect 683 2254 692 2263
rect 797 2254 806 2263
rect 911 2254 920 2263
rect 1025 2254 1034 2263
rect 1139 2254 1148 2263
rect 1253 2254 1262 2263
rect 1832 1795 1837 1800
rect 2332 1795 2337 1800
rect 3002 1603 3007 1608
rect 1083 1563 1092 1572
rect 75 903 84 912
rect 105 603 112 612
<< metal3 >>
rect 75 3012 84 3353
rect 75 2662 84 3003
rect 1640 2993 1645 3309
rect 1679 3133 1684 3291
rect 2597 3285 2600 3291
rect 1679 3128 1714 3133
rect 1679 3111 1684 3128
rect 1665 3106 1684 3111
rect 1717 3094 1722 3107
rect 1668 3089 1722 3094
rect 1738 3080 1743 3128
rect 1656 3075 1743 3080
rect 1640 2988 1661 2993
rect 1587 2967 1705 2972
rect 1568 2962 1577 2965
rect 1568 2953 2416 2962
rect 1587 2902 2317 2911
rect 2308 2892 2317 2902
rect 2308 2883 2367 2892
rect 2407 2859 2416 2953
rect 1336 2791 1339 2796
rect 75 2312 84 2653
rect 75 1962 84 2303
rect 2591 2242 2600 3285
rect 1863 2232 2352 2242
rect 2363 2232 2600 2242
rect 75 1612 84 1953
rect 75 1262 84 1603
rect 411 2196 2699 2205
rect 411 1601 420 2196
rect 453 2195 483 2196
rect 532 2178 2717 2187
rect 532 1576 541 2178
rect 885 2160 2735 2169
rect 885 1684 894 2160
rect 917 2142 2763 2151
rect 917 1684 926 2142
rect 951 2124 2781 2133
rect 951 1684 960 2124
rect 1057 2106 2799 2115
rect 1057 1706 1066 2106
rect 1083 2088 2817 2097
rect 986 1684 991 1689
rect 986 1653 991 1662
rect 715 1621 720 1626
rect 777 1621 782 1626
rect 936 1574 941 1653
rect 1083 1572 1092 2088
rect 1205 2070 2845 2079
rect 1205 1815 1214 2070
rect 1205 1634 1214 1810
rect 1225 2052 2863 2061
rect 1205 1625 1207 1634
rect 1225 1625 1234 2052
rect 1403 2034 2881 2043
rect 1403 1625 1412 2034
rect 1488 2016 2899 2025
rect 1488 1741 1497 2016
rect 1512 1998 2927 2007
rect 1512 1625 1521 1998
rect 1356 1616 1388 1621
rect 1403 1616 1436 1625
rect 1461 1616 1521 1625
rect 1534 1980 2945 1989
rect 1534 1616 1543 1980
rect 1641 1962 2963 1971
rect 1564 1616 1602 1621
rect 1641 1616 1650 1962
rect 1671 1616 1709 1621
rect 1748 1616 1757 1962
rect 1830 1944 2981 1953
rect 1830 1800 1842 1944
rect 1875 1926 3009 1935
rect 1875 1620 1884 1926
rect 1948 1908 3027 1917
rect 1429 1612 1434 1616
rect 1463 1612 1468 1616
rect 1536 1612 1541 1616
rect 1570 1612 1575 1616
rect 1597 1612 1602 1616
rect 1643 1612 1648 1616
rect 1677 1612 1682 1616
rect 1704 1611 1709 1616
rect 1750 1612 1755 1616
rect 1877 1615 1882 1620
rect 1948 1615 1957 1908
rect 2200 1890 3045 1899
rect 2200 1622 2209 1890
rect 2330 1872 3063 1881
rect 2330 1800 2342 1872
rect 2448 1854 3091 1863
rect 1950 1612 1955 1615
rect 2375 1620 2384 1746
rect 2200 1608 2209 1613
rect 2377 1612 2382 1620
rect 2448 1615 2457 1854
rect 2482 1836 3109 1845
rect 2482 1616 2491 1836
rect 2555 1818 3127 1827
rect 2555 1616 2564 1818
rect 2675 1800 3145 1809
rect 2675 1616 2684 1800
rect 2748 1782 3173 1791
rect 3218 1782 3396 1791
rect 2748 1616 2757 1782
rect 3124 1764 3189 1773
rect 3198 1764 3258 1773
rect 2450 1612 2455 1615
rect 2484 1612 2489 1616
rect 2557 1612 2562 1616
rect 2677 1612 2682 1616
rect 2750 1612 2755 1616
rect 3124 1608 3133 1764
rect 3248 1608 3258 1764
rect 411 1568 416 1571
rect 536 1568 541 1571
rect 859 1561 864 1566
rect 1066 1561 1071 1566
rect 1327 1564 1332 1569
rect 2202 1568 2207 1574
rect 3002 1570 3007 1574
rect 3126 1571 3131 1575
rect 3250 1569 3255 1573
rect 75 912 84 1253
rect 84 903 121 912
rect 3386 905 3396 1782
rect 112 612 121 903
rect 112 603 325 612
rect 311 222 325 603
rect 3385 435 3396 905
rect 3385 222 3395 435
rect 311 209 3395 222
rect 311 208 325 209
<< m234contact >>
rect 1006 3585 1015 3594
rect 1658 3282 1668 3291
rect 1360 2896 1369 2905
rect 2475 2896 2485 2905
rect 1360 2832 1369 2841
rect 2451 2832 2460 2841
rect 1674 2791 1679 2796
rect 2344 2777 2353 2786
rect 1360 2768 1369 2777
rect 1360 2704 1369 2713
rect 2308 2704 2317 2713
rect 3557 2726 3566 2735
rect 3557 2376 3566 2385
rect 859 1606 864 1611
rect 878 1592 883 1597
rect 1296 1820 1301 1825
rect 1309 1810 1314 1815
rect 3557 2026 3566 2035
rect 1465 1635 1470 1640
rect 1343 1616 1352 1625
rect 1866 1615 1871 1620
rect 1452 1605 1457 1610
rect 1490 1605 1495 1610
rect 2473 1607 2478 1612
rect 3186 1572 3194 1580
rect 478 1546 483 1551
rect 878 1416 883 1421
rect 3186 1396 3194 1404
rect 478 1370 483 1375
rect 878 1240 883 1245
rect 3186 1220 3194 1228
rect 478 1194 483 1199
rect 878 1064 883 1069
rect 3186 1044 3194 1052
rect 478 1018 483 1023
rect 3557 1676 3566 1685
rect 3557 1326 3566 1335
rect 3557 976 3566 985
rect 878 888 883 893
rect 3186 868 3194 876
rect 478 842 483 847
rect 878 712 883 717
rect 3186 692 3194 700
rect 478 666 483 671
rect 878 536 883 541
rect 3186 516 3194 524
rect 478 490 483 495
rect 3557 626 3566 635
rect 878 360 883 365
rect 3186 340 3194 348
rect 478 314 483 319
rect 3557 276 3566 285
<< m4contact >>
rect 1640 3309 1645 3314
rect 1679 3291 1684 3296
rect 2591 3291 2600 3300
rect 2642 3291 2651 3300
rect 1413 2955 1422 2964
rect 1531 2955 1540 2964
rect 1339 2791 1344 2796
rect 1852 2232 1863 2242
rect 2352 2232 2363 2242
rect 936 1653 941 1658
rect 981 1653 986 1658
rect 1205 1810 1214 1815
rect 1207 1625 1216 1634
rect 1225 1616 1234 1625
rect 1857 1738 1862 1743
rect 2357 1738 2362 1743
rect 2200 1613 2209 1622
rect 2511 1607 2516 1612
rect 469 1506 474 1511
rect 469 1330 474 1335
rect 469 1154 474 1159
rect 469 978 474 983
rect 469 802 474 807
rect 469 626 474 631
rect 469 450 474 455
rect 469 274 474 279
<< metal4 >>
rect 1006 3320 1015 3585
rect 1006 3319 1330 3320
rect 1006 3318 1454 3319
rect 1006 3314 2651 3318
rect 1006 3311 1640 3314
rect 1227 3310 1640 3311
rect 1413 3309 1640 3310
rect 1645 3309 2651 3314
rect 1413 2964 1422 3309
rect 2642 3300 2651 3309
rect 1531 3296 2591 3300
rect 1531 3291 1679 3296
rect 1684 3291 2591 3296
rect 1531 2964 1540 3291
rect 1369 2896 2475 2905
rect 1369 2832 2451 2841
rect 1344 2791 1674 2796
rect 1369 2768 2353 2777
rect 3280 2735 3529 2744
rect 3280 2726 3557 2735
rect 3280 2721 3529 2726
rect 1369 2704 2308 2713
rect 3280 2679 3308 2721
rect 1301 1820 1470 1825
rect 1214 1810 1309 1815
rect 941 1653 981 1658
rect 1465 1640 1470 1820
rect 1852 1743 1863 2232
rect 2352 1743 2363 2232
rect 1852 1738 1857 1743
rect 1862 1738 1863 1743
rect 3182 1702 3199 1705
rect 3279 1702 3308 2679
rect 3181 1685 3308 1702
rect 3334 2387 3515 2388
rect 3334 2385 3516 2387
rect 3334 2376 3557 2385
rect 3334 2372 3516 2376
rect 3181 1684 3302 1685
rect 1234 1616 1343 1625
rect 1871 1613 2200 1622
rect 1457 1605 1490 1610
rect 2478 1607 2511 1612
rect 3182 1580 3199 1684
rect 3334 1405 3358 2372
rect 3194 1396 3358 1405
rect 3334 1394 3358 1396
rect 3377 2035 3397 2036
rect 3377 2026 3557 2035
rect 3377 2022 3531 2026
rect 3377 1229 3397 2022
rect 3194 1220 3397 1229
rect 3377 1216 3397 1220
rect 3422 1687 3438 1688
rect 3422 1686 3439 1687
rect 3422 1685 3522 1686
rect 3422 1676 3557 1685
rect 3422 1675 3522 1676
rect 3422 1053 3439 1675
rect 3194 1044 3439 1053
rect 3422 1043 3439 1044
rect 3465 1326 3557 1335
rect 3465 877 3479 1326
rect 3506 985 3517 986
rect 3506 976 3557 985
rect 3506 877 3517 976
rect 3194 868 3479 877
rect 3505 868 3517 877
rect 3465 866 3479 868
rect 3506 701 3517 868
rect 3194 692 3517 701
rect 3506 626 3557 635
rect 3506 525 3517 626
rect 3194 516 3517 525
rect 3186 348 3517 349
rect 3194 340 3517 348
rect 3506 285 3517 340
rect 3506 277 3557 285
rect 3507 276 3557 277
<< m345contact >>
rect 455 2244 464 2254
rect 569 2244 578 2253
rect 683 2245 692 2254
rect 797 2245 806 2254
rect 911 2245 920 2254
rect 1025 2245 1034 2254
rect 1139 2245 1148 2254
rect 1253 2245 1262 2254
rect 3318 1548 3326 1557
rect 3318 1372 3326 1381
rect 3318 1196 3326 1205
rect 3318 1020 3326 1029
rect 3318 844 3326 853
rect 3318 668 3326 677
rect 3318 492 3326 501
rect 3318 316 3326 325
rect 607 102 616 110
rect 957 102 966 110
rect 1307 102 1316 110
rect 1657 102 1666 110
rect 2007 102 2016 110
rect 2357 102 2366 110
rect 2707 102 2716 110
rect 3057 102 3066 110
<< m5contact >>
rect 476 1551 485 1560
rect 476 1375 485 1384
rect 476 1199 485 1208
rect 476 1023 485 1032
rect 476 847 485 856
rect 476 671 485 680
rect 476 495 485 504
rect 476 319 485 328
<< metal5 >>
rect 455 1560 464 2244
rect 455 1551 476 1560
rect 569 1384 578 2244
rect 485 1375 579 1384
rect 683 1208 692 2245
rect 485 1199 692 1208
rect 797 1032 806 2245
rect 485 1023 806 1032
rect 911 856 920 2245
rect 485 847 920 856
rect 1025 680 1034 2245
rect 485 671 1034 680
rect 1139 504 1148 2245
rect 485 495 1148 504
rect 1139 494 1148 495
rect 1253 328 1262 2245
rect 1519 1563 3333 1564
rect 1333 1557 3333 1563
rect 1333 1548 3318 1557
rect 3326 1548 3333 1557
rect 1333 1544 3333 1548
rect 1332 1539 3333 1544
rect 1332 1537 1632 1539
rect 1332 1195 1352 1537
rect 1519 1387 3333 1389
rect 1436 1383 3333 1387
rect 1429 1381 3333 1383
rect 1429 1372 3318 1381
rect 3326 1372 3333 1381
rect 1429 1364 3333 1372
rect 1429 1358 1565 1364
rect 485 319 1262 328
rect 1335 304 1349 1195
rect 1429 1133 1444 1358
rect 1516 1206 1535 1209
rect 1513 1205 3327 1206
rect 1513 1196 3318 1205
rect 3326 1196 3327 1205
rect 1513 1181 3327 1196
rect 1428 1116 1444 1133
rect 1335 246 1351 304
rect 1428 263 1442 1116
rect 1516 1001 1535 1181
rect 1653 1029 3343 1038
rect 1653 1020 3318 1029
rect 3326 1020 3343 1029
rect 1653 1001 3343 1020
rect 604 226 1355 246
rect 604 225 1092 226
rect 607 110 620 225
rect 1424 182 1444 263
rect 958 164 1446 182
rect 616 102 620 110
rect 957 161 1446 164
rect 957 110 966 161
rect 1307 137 1316 139
rect 1517 137 1531 1001
rect 1307 118 1531 137
rect 1657 998 1690 1001
rect 1307 117 1503 118
rect 1307 110 1316 117
rect 1657 110 1671 998
rect 2001 853 3334 856
rect 2001 844 3318 853
rect 3326 844 3334 853
rect 2001 842 3334 844
rect 1666 102 1671 110
rect 2007 110 2029 842
rect 2354 677 3328 687
rect 2354 668 3318 677
rect 3326 668 3328 677
rect 2354 663 3328 668
rect 2016 102 2029 110
rect 2357 110 2368 663
rect 2709 501 3328 506
rect 2709 492 3318 501
rect 3326 492 3328 501
rect 2709 485 3328 492
rect 2366 102 2368 110
rect 2707 484 3328 485
rect 2707 110 2717 484
rect 3230 316 3318 325
rect 3230 114 3244 316
rect 2716 102 2717 110
rect 3057 110 3244 114
rect 3066 102 3244 110
use inv2  inv2_0
timestamp 1765746878
transform -1 0 95 0 -1 618
box -10 -13 20 40
use datapath  datapath_0
timestamp 1765789580
transform 1 0 431 0 1 -264
box -81 532 2885 2021
use latch_one  latch_one_0
timestamp 1765002978
transform 0 -1 1796 -1 0 1779
box -11 -67 48 -12
use latch_one  latch_one_1
timestamp 1765002978
transform 0 -1 2296 -1 0 1779
box -11 -67 48 -12
use 2and  2and_0
timestamp 1765747547
transform -1 0 1396 0 1 1729
box 68 29 138 82
use control  control_0
timestamp 1765789580
transform -1 0 1314 0 -1 3151
box -317 -140 974 447
use rom  rom_0
timestamp 1765759847
transform 1 0 2676 0 1 3129
box -350 -907 584 162
use 4nor  4nor_0
timestamp 1765673320
transform 0 1 1666 -1 0 3295
box 72 -6 132 47
use inv  inv_0
timestamp 1765001281
transform 0 1 1673 -1 0 3243
box -10 -13 20 40
use inv  inv_1
timestamp 1765001281
transform 1 0 1724 0 1 3117
box -10 -13 20 40
use 2and  2and_1
timestamp 1765747547
transform 0 1 1631 -1 0 3054
box 68 29 138 82
use staticizer_one  staticizer_one_0
timestamp 1765746506
transform 0 1 1717 -1 0 3158
box 54 -61 113 -1
use latch_one  latch_one_2
timestamp 1765002978
transform 0 1 1726 -1 0 3152
box -11 -67 48 -12
use latch_one  latch_one_3
timestamp 1765002978
transform 0 1 1725 -1 0 3034
box -11 -67 48 -12
use 0names  0names_0
timestamp 1765780088
transform 1 0 1777 0 1 2432
box -128 -44 222 94
use ring  ring_0
timestamp 1765052771
transform 1 0 179 0 1 3594
box -207 -3603 3499 111
<< labels >>
rlabel metal1 351 1209 356 1214 3 data_out2
rlabel metal1 351 1033 356 1038 3 data_out3
rlabel metal1 351 857 356 862 3 data_out4
rlabel metal1 351 681 356 686 3 data_out5
rlabel metal1 351 505 356 510 3 data_out6
rlabel metal1 351 329 356 334 3 data_out7
rlabel m234contact 478 314 483 319 1 data_in7
rlabel m234contact 478 490 483 495 1 data_in6
rlabel m234contact 478 666 483 671 1 data_in5
rlabel m234contact 478 842 483 847 1 data_in4
rlabel m234contact 478 1018 483 1023 1 data_in3
rlabel m234contact 478 1194 483 1199 1 data_in2
rlabel m234contact 478 1370 483 1375 1 data_in1
rlabel metal2 3209 2045 3218 2054 1 r_-w
rlabel metal1 3254 1359 3259 1364 1 addr_out9
rlabel metal1 3254 1535 3259 1540 1 addr_out8
rlabel metal1 3254 1183 3259 1188 1 addr_out10
rlabel metal1 3254 1007 3259 1012 1 addr_out11
rlabel metal1 3254 831 3259 836 1 addr_out12
rlabel metal1 3254 655 3259 660 1 addr_out13
rlabel metal1 3254 479 3259 484 1 addr_out14
rlabel metal1 3254 303 3259 308 1 addr_out15
rlabel metal1 3130 1536 3135 1540 1 addr_out0
rlabel metal1 3130 1360 3135 1364 1 addr_out1
rlabel metal1 3130 1184 3135 1188 1 addr_out2
rlabel metal1 3130 1008 3135 1012 1 addr_out3
rlabel metal1 3130 832 3135 836 1 addr_out4
rlabel metal1 3130 656 3135 660 1 addr_out5
rlabel metal1 3130 480 3135 484 1 addr_out6
rlabel metal1 3130 304 3135 308 1 addr_out7
rlabel metal1 2360 2546 2365 2551 1 s3
rlabel metal1 2380 2595 2385 2600 1 s2
rlabel metal1 2460 3134 2465 3139 1 s1
rlabel metal1 2470 3087 2475 3092 1 s0
rlabel metal3 411 1568 416 1571 1 rd_dataout
rlabel metal3 536 1568 541 1571 1 ld_datain
rlabel metal3 715 1621 720 1626 1 os_u
rlabel metal3 777 1621 782 1626 1 os_s
rlabel metal3 859 1561 864 1566 1 ros
rlabel metal3 887 1684 892 1689 1 fb_g3
rlabel metal3 919 1684 924 1689 1 fb_g2
rlabel metal3 953 1684 958 1689 1 fb_g1
rlabel metal3 986 1684 991 1689 1 fb_g0
rlabel metal3 1066 1561 1071 1566 1 rfb
rlabel m123contact 1087 1565 1092 1570 1 as_sub
rlabel metal1 1273 1634 1278 1639 1 as_cin
rlabel m234contact 1345 1616 1350 1621 1 A_r0
rlabel metal3 1356 1616 1361 1621 1 A_r1
rlabel metal3 1327 1564 1332 1569 1 ras
rlabel m234contact 878 1592 883 1597 1 ry0
rlabel m234contact 878 1416 883 1421 1 ry1
rlabel m234contact 878 1240 883 1245 1 ry2
rlabel m234contact 878 1064 883 1069 1 ry3
rlabel m234contact 878 888 883 893 1 ry4
rlabel m234contact 878 712 883 717 1 ry5
rlabel m234contact 878 536 883 541 1 ry6
rlabel m234contact 878 360 883 365 1 ry7
rlabel m4contact 469 1506 474 1511 1 rx0
rlabel m4contact 469 1330 474 1335 1 rx1
rlabel m4contact 469 1154 474 1159 1 rx2
rlabel m4contact 469 978 474 983 1 rx3
rlabel m4contact 469 802 474 807 1 rx4
rlabel m4contact 469 626 474 631 1 rx5
rlabel m4contact 469 450 474 455 1 rx6
rlabel m4contact 469 274 474 279 1 rx7
rlabel m2contact 1959 1523 1964 1526 1 rx_PCL0
rlabel m2contact 1959 1347 1964 1350 1 rx_PCL1
rlabel m2contact 1959 1171 1964 1174 1 rx_PCL2
rlabel m2contact 1959 995 1964 998 1 rx_PCL3
rlabel m2contact 1959 819 1964 822 1 rx_PCL4
rlabel m2contact 1959 643 1964 646 1 rx_PCL5
rlabel m2contact 1959 467 1964 470 1 rx_PCL6
rlabel m2contact 1959 291 1964 294 1 rx_PCL7
rlabel metal3 1429 1612 1434 1616 1 A_w
rlabel metal2 1452 1612 1457 1616 1 DB_r0
rlabel metal3 1463 1612 1468 1616 1 DB_r1
rlabel metal3 1536 1612 1541 1616 1 DB_w
rlabel metal2 1559 1612 1564 1616 1 X_r0
rlabel metal3 1570 1612 1575 1616 1 X_r1
rlabel metal3 1643 1612 1648 1616 1 X_w
rlabel metal2 1666 1612 1671 1616 1 Y_r0
rlabel metal3 1677 1612 1682 1616 1 Y_r1
rlabel metal3 1750 1612 1755 1616 1 Y_w
rlabel metal3 1876 1622 1881 1627 1 PCL_r1
rlabel metal2 1866 1612 1871 1615 1 PCL_r0
rlabel metal3 1950 1612 1955 1615 1 PCL_w
rlabel metal3 2202 1571 2207 1574 1 rPCplus1L
rlabel metal2 2366 1612 2371 1615 1 PCH_r0
rlabel metal3 2377 1612 2382 1615 1 PCH_r1
rlabel metal3 2450 1612 2455 1615 1 PCH_w
rlabel metal2 2473 1612 2478 1616 1 ABL_r0
rlabel metal3 2484 1612 2489 1616 1 ABL_r1
rlabel metal3 2557 1612 2562 1616 1 ABL_w
rlabel metal1 2635 1732 2640 1736 1 ABH_w_sel
rlabel metal2 2666 1612 2671 1616 1 ABH_r0
rlabel metal3 2677 1612 2682 1616 1 ABH_r1
rlabel metal3 2750 1612 2755 1616 1 ABH_w
rlabel metal3 3002 1570 3007 1574 1 rPCplus1H
rlabel metal3 3126 1572 3131 1575 1 rd_addrL
rlabel metal3 3250 1570 3255 1573 1 rd_addrH
rlabel metal1 2335 1729 2339 1732 1 PCH_w_sel
rlabel metal1 1835 1725 1840 1732 1 PCL_w_sel
rlabel metal3 1491 1741 1496 1746 1 Cflag_w
rlabel m2contact 1489 1638 1494 1643 1 Cflag
rlabel space 177 3682 319 3696 1 Vdd!
rlabel space 632 3688 640 3700 1 phi0
rlabel space 982 3690 990 3702 1 phi1
rlabel space 1332 3688 1340 3705 1 reset
rlabel space -29 3452 -17 3460 1 r-w_
rlabel space -29 3102 -17 3110 1 d0
rlabel space -29 2752 -17 2760 1 d1
rlabel space -29 2402 -17 2410 1 d2
rlabel space -29 2052 -17 2060 1 d3
rlabel space -29 1702 -17 1710 1 d4
rlabel space -29 1352 -18 1360 1 d5
rlabel space -29 1002 -17 1010 1 d6
rlabel space -29 652 -17 660 1 d7
rlabel space -28 198 -14 340 1 GND!
rlabel space 558 -9 566 3 1 a15
rlabel space 908 -9 916 3 1 a14
rlabel space 1258 -9 1266 3 1 a13
rlabel space 1608 -9 1616 3 1 a12
rlabel space 1958 -9 1966 3 1 a11
rlabel space 2308 -9 2316 3 1 a10
rlabel space 2658 -9 2666 3 1 a9
rlabel space 3008 -9 3016 3 1 a8
rlabel space 3328 -8 3470 6 1 Vdd!
rlabel space 3665 228 3677 236 1 a7
rlabel space 3665 578 3677 586 1 a6
rlabel space 3665 928 3677 936 1 a5
rlabel space 3665 1278 3677 1286 1 a4
rlabel space 3665 1628 3677 1636 1 a3
rlabel space 3665 1978 3677 1986 1 a2
rlabel space 3665 2328 3677 2336 1 a1
rlabel space 3665 2678 3677 2686 1 a0
rlabel space 3662 3348 3676 3490 1 GND!
rlabel m234contact 478 1546 483 1551 1 data_in0
rlabel metal1 1331 3254 1336 3259 1 rst
rlabel metal2 528 2800 533 2803 1 IR0
rlabel metal2 642 2800 647 2803 1 IR1
rlabel metal2 756 2799 761 2802 1 IR2
rlabel metal2 870 2800 875 2803 1 IR3
rlabel metal2 984 2800 989 2803 1 IR4
rlabel metal2 1098 2785 1103 2788 1 IR5
rlabel metal2 1212 2799 1217 2802 1 IR6
rlabel metal2 1326 2799 1331 2802 1 IR7
rlabel metal2 749 3259 754 3262 1 s0'
rlabel metal2 603 3259 608 3262 1 s1'
rlabel metal2 448 3259 453 3262 1 s2'
rlabel metal1 1474 2925 1479 2930 1 s0_int
rlabel metal1 1474 2861 1479 2866 1 s1_int
rlabel metal1 1474 2797 1479 2802 1 s2_int
rlabel metal1 1474 2733 1479 2738 1 s3_int
rlabel metal2 340 3259 345 3262 1 s3'
rlabel polycontact 1685 3162 1690 3167 1 IR_w_next
rlabel m4contact 1339 2791 1344 2796 1 IR_w
rlabel polycontact 1684 3102 1689 3107 1 IR_w_int
rlabel polycontact 1681 2981 1686 2986 1 IR_w_latched
rlabel metal1 3575 676 3582 685 7 ring_0/pad_6[8]/oe
rlabel metal1 3575 1026 3582 1035 7 ring_0/pad_6[8]/oe
rlabel metal1 3575 1376 3582 1385 7 ring_0/pad_6[8]/oe
rlabel metal1 3575 1726 3582 1735 7 ring_0/pad_6[8]/oe
rlabel metal1 3575 2076 3582 2085 7 ring_0/pad_6[8]/oe
rlabel metal1 3575 2426 3582 2435 7 ring_0/pad_6[8]/oe
rlabel metal1 3575 2776 3582 2785 7 ring_0/pad_6[8]/oe
<< end >>
