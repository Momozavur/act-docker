magic
tech scmos
timestamp 1765747812
<< nwell >>
rect 72 52 120 81
<< pwell >>
rect 72 28 120 51
<< ntransistor >>
rect 85 40 87 45
rect 95 40 97 45
rect 106 40 108 45
<< ptransistor >>
rect 85 58 87 69
rect 95 58 97 69
rect 106 58 108 69
<< ndiffusion >>
rect 83 40 85 45
rect 87 40 89 45
rect 94 40 95 45
rect 97 40 99 45
rect 104 40 106 45
rect 108 40 109 45
<< pdiffusion >>
rect 83 58 85 69
rect 87 58 95 69
rect 97 58 106 69
rect 108 58 109 69
<< ndcontact >>
rect 78 40 83 45
rect 89 40 94 45
rect 99 40 104 45
rect 109 40 114 45
<< pdcontact >>
rect 78 58 83 69
rect 109 58 114 69
<< psubstratepcontact >>
rect 99 31 104 36
<< nsubstratencontact >>
rect 99 73 104 78
<< polysilicon >>
rect 85 69 87 72
rect 95 69 97 72
rect 106 69 108 72
rect 85 45 87 58
rect 95 45 97 58
rect 106 45 108 58
rect 85 37 87 40
rect 95 37 97 40
rect 106 37 108 40
<< metal1 >>
rect 78 73 99 78
rect 104 73 120 78
rect 78 69 83 73
rect 109 54 114 58
rect 89 49 120 54
rect 89 45 94 49
rect 109 45 114 49
rect 78 36 83 40
rect 99 36 104 40
rect 78 31 99 36
rect 104 31 120 36
<< labels >>
rlabel polysilicon 85 70 87 72 1 a
rlabel polysilicon 95 70 97 72 1 b
rlabel metal1 115 49 120 54 7 out
rlabel metal1 115 31 120 36 7 GND!
rlabel polysilicon 106 70 108 72 1 c
rlabel metal1 115 73 120 78 7 Vdd!
<< end >>
